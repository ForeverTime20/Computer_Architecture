��` t i m e s c a l e   1 n s / 1 0 0 p s  
 / / c o r r e c t   r e a d   r e s u l t :  
 / /   0 0 0 0 0 0 2 9   0 0 0 0 0 0 0 6   0 0 0 0 0 0 1 0   0 0 0 0 0 0 1 2   0 0 0 0 0 0 0 e   0 0 0 0 0 0 0 4   0 0 0 0 0 0 1 0   0 0 0 0 0 0 1 7   0 0 0 0 0 0 0 9   0 0 0 0 0 0 0 b   0 0 0 0 0 0 1 e   0 0 0 0 0 0 2 6   0 0 0 0 0 0 0 4   0 0 0 0 0 0 3 e   0 0 0 0 0 0 0 2   0 0 0 0 0 0 1 4  
  
 m o d u l e   c a c h e _ t b ( ) ;  
  
 ` d e f i n e   D A T A _ C O U N T   ( 1 6 )  
 ` d e f i n e   R D W R _ C O U N T   ( 6 * ` D A T A _ C O U N T )  
  
 r e g   w r _ c y c l e                       [ ` R D W R _ C O U N T ] ;  
 r e g   r d _ c y c l e                       [ ` R D W R _ C O U N T ] ;  
 r e g   [ 3 1 : 0 ]   a d d r _ r o m         [ ` R D W R _ C O U N T ] ;  
 r e g   [ 3 1 : 0 ]   w r _ d a t a _ r o m   [ ` R D W R _ C O U N T ] ;  
 r e g   [ 3 1 : 0 ]   v a l i d a t i o n _ d a t a   [ ` D A T A _ C O U N T ] ;  
  
 i n i t i a l   b e g i n  
         / /   1 6   s e q u e n c e   w r i t e   c y c l e s  
         r d _ c y c l e [         0 ]   =   1 ' b 0 ;     w r _ c y c l e [         0 ]   =   1 ' b 1 ;     a d d r _ r o m [         0 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [         0 ] = ' h 0 0 0 0 0 0 1 c ;  
         r d _ c y c l e [         1 ]   =   1 ' b 0 ;     w r _ c y c l e [         1 ]   =   1 ' b 1 ;     a d d r _ r o m [         1 ] = ' h 0 0 0 0 0 0 0 4 ;     w r _ d a t a _ r o m [         1 ] = ' h 0 0 0 0 0 0 1 b ;  
         r d _ c y c l e [         2 ]   =   1 ' b 0 ;     w r _ c y c l e [         2 ]   =   1 ' b 1 ;     a d d r _ r o m [         2 ] = ' h 0 0 0 0 0 0 0 8 ;     w r _ d a t a _ r o m [         2 ] = ' h 0 0 0 0 0 0 1 8 ;  
         r d _ c y c l e [         3 ]   =   1 ' b 0 ;     w r _ c y c l e [         3 ]   =   1 ' b 1 ;     a d d r _ r o m [         3 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [         3 ] = ' h 0 0 0 0 0 0 2 b ;  
         r d _ c y c l e [         4 ]   =   1 ' b 0 ;     w r _ c y c l e [         4 ]   =   1 ' b 1 ;     a d d r _ r o m [         4 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [         4 ] = ' h 0 0 0 0 0 0 2 8 ;  
         r d _ c y c l e [         5 ]   =   1 ' b 0 ;     w r _ c y c l e [         5 ]   =   1 ' b 1 ;     a d d r _ r o m [         5 ] = ' h 0 0 0 0 0 0 1 4 ;     w r _ d a t a _ r o m [         5 ] = ' h 0 0 0 0 0 0 1 5 ;  
         r d _ c y c l e [         6 ]   =   1 ' b 0 ;     w r _ c y c l e [         6 ]   =   1 ' b 1 ;     a d d r _ r o m [         6 ] = ' h 0 0 0 0 0 0 1 8 ;     w r _ d a t a _ r o m [         6 ] = ' h 0 0 0 0 0 0 1 6 ;  
         r d _ c y c l e [         7 ]   =   1 ' b 0 ;     w r _ c y c l e [         7 ]   =   1 ' b 1 ;     a d d r _ r o m [         7 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [         7 ] = ' h 0 0 0 0 0 0 1 9 ;  
         r d _ c y c l e [         8 ]   =   1 ' b 0 ;     w r _ c y c l e [         8 ]   =   1 ' b 1 ;     a d d r _ r o m [         8 ] = ' h 0 0 0 0 0 0 2 0 ;     w r _ d a t a _ r o m [         8 ] = ' h 0 0 0 0 0 0 4 0 ;  
         r d _ c y c l e [         9 ]   =   1 ' b 0 ;     w r _ c y c l e [         9 ]   =   1 ' b 1 ;     a d d r _ r o m [         9 ] = ' h 0 0 0 0 0 0 2 4 ;     w r _ d a t a _ r o m [         9 ] = ' h 0 0 0 0 0 0 3 f ;  
         r d _ c y c l e [       1 0 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 0 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 0 ] = ' h 0 0 0 0 0 0 2 8 ;     w r _ d a t a _ r o m [       1 0 ] = ' h 0 0 0 0 0 0 1 e ;  
         r d _ c y c l e [       1 1 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 1 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 1 ] = ' h 0 0 0 0 0 0 2 c ;     w r _ d a t a _ r o m [       1 1 ] = ' h 0 0 0 0 0 0 3 2 ;  
         r d _ c y c l e [       1 2 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 2 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 2 ] = ' h 0 0 0 0 0 0 3 0 ;     w r _ d a t a _ r o m [       1 2 ] = ' h 0 0 0 0 0 0 3 3 ;  
         r d _ c y c l e [       1 3 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 3 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 3 ] = ' h 0 0 0 0 0 0 3 4 ;     w r _ d a t a _ r o m [       1 3 ] = ' h 0 0 0 0 0 0 3 e ;  
         r d _ c y c l e [       1 4 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 4 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 4 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       1 4 ] = ' h 0 0 0 0 0 0 1 9 ;  
         r d _ c y c l e [       1 5 ]   =   1 ' b 0 ;     w r _ c y c l e [       1 5 ]   =   1 ' b 1 ;     a d d r _ r o m [       1 5 ] = ' h 0 0 0 0 0 0 3 c ;     w r _ d a t a _ r o m [       1 5 ] = ' h 0 0 0 0 0 0 1 4 ;  
         / /   4 8   r a n d o m   r e a d   a n d   w r i t e   c y c l e s  
         r d _ c y c l e [       1 6 ]   =   1 ' b 1 ;     w r _ c y c l e [       1 6 ]   =   1 ' b 0 ;     a d d r _ r o m [       1 6 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       1 6 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       1 7 ]   =   1 ' b 1 ;     w r _ c y c l e [       1 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       1 7 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       1 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       1 8 ]   =   1 ' b 1 ;     w r _ c y c l e [       1 8 ]   =   1 ' b 0 ;     a d d r _ r o m [       1 8 ] = ' h 0 0 0 0 0 0 0 8 ;     w r _ d a t a _ r o m [       1 8 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       1 9 ]   =   1 ' b 1 ;     w r _ c y c l e [       1 9 ]   =   1 ' b 0 ;     a d d r _ r o m [       1 9 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [       1 9 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 0 ]   =   1 ' b 0 ;     w r _ c y c l e [       2 0 ]   =   1 ' b 1 ;     a d d r _ r o m [       2 0 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       2 0 ] = ' h 0 0 0 0 0 0 1 e ;  
         r d _ c y c l e [       2 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       2 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       2 1 ] = ' h 0 0 0 0 0 0 1 8 ;     w r _ d a t a _ r o m [       2 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 2 ]   =   1 ' b 1 ;     w r _ c y c l e [       2 2 ]   =   1 ' b 0 ;     a d d r _ r o m [       2 2 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [       2 2 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       2 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       2 3 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       2 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 4 ]   =   1 ' b 0 ;     w r _ c y c l e [       2 4 ]   =   1 ' b 1 ;     a d d r _ r o m [       2 4 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       2 4 ] = ' h 0 0 0 0 0 0 3 5 ;  
         r d _ c y c l e [       2 5 ]   =   1 ' b 1 ;     w r _ c y c l e [       2 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       2 5 ] = ' h 0 0 0 0 0 0 3 c ;     w r _ d a t a _ r o m [       2 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 6 ]   =   1 ' b 0 ;     w r _ c y c l e [       2 6 ]   =   1 ' b 1 ;     a d d r _ r o m [       2 6 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       2 6 ] = ' h 0 0 0 0 0 0 0 e ;  
         r d _ c y c l e [       2 7 ]   =   1 ' b 1 ;     w r _ c y c l e [       2 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       2 7 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       2 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       2 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       2 8 ]   =   1 ' b 1 ;     a d d r _ r o m [       2 8 ] = ' h 0 0 0 0 0 0 2 c ;     w r _ d a t a _ r o m [       2 8 ] = ' h 0 0 0 0 0 0 2 6 ;  
         r d _ c y c l e [       2 9 ]   =   1 ' b 0 ;     w r _ c y c l e [       2 9 ]   =   1 ' b 1 ;     a d d r _ r o m [       2 9 ] = ' h 0 0 0 0 0 0 1 4 ;     w r _ d a t a _ r o m [       2 9 ] = ' h 0 0 0 0 0 0 0 4 ;  
         r d _ c y c l e [       3 0 ]   =   1 ' b 1 ;     w r _ c y c l e [       3 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       3 0 ] = ' h 0 0 0 0 0 0 3 0 ;     w r _ d a t a _ r o m [       3 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       3 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       3 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       3 1 ] = ' h 0 0 0 0 0 0 3 4 ;     w r _ d a t a _ r o m [       3 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       3 2 ]   =   1 ' b 0 ;     w r _ c y c l e [       3 2 ]   =   1 ' b 1 ;     a d d r _ r o m [       3 2 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [       3 2 ] = ' h 0 0 0 0 0 0 1 d ;  
         r d _ c y c l e [       3 3 ]   =   1 ' b 0 ;     w r _ c y c l e [       3 3 ]   =   1 ' b 1 ;     a d d r _ r o m [       3 3 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       3 3 ] = ' h 0 0 0 0 0 0 1 6 ;  
         r d _ c y c l e [       3 4 ]   =   1 ' b 1 ;     w r _ c y c l e [       3 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       3 4 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       3 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       3 5 ]   =   1 ' b 1 ;     w r _ c y c l e [       3 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       3 5 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       3 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       3 6 ]   =   1 ' b 0 ;     w r _ c y c l e [       3 6 ]   =   1 ' b 1 ;     a d d r _ r o m [       3 6 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [       3 6 ] = ' h 0 0 0 0 0 0 1 2 ;  
         r d _ c y c l e [       3 7 ]   =   1 ' b 1 ;     w r _ c y c l e [       3 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       3 7 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [       3 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       3 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       3 8 ]   =   1 ' b 1 ;     a d d r _ r o m [       3 8 ] = ' h 0 0 0 0 0 0 1 8 ;     w r _ d a t a _ r o m [       3 8 ] = ' h 0 0 0 0 0 0 1 0 ;  
         r d _ c y c l e [       3 9 ]   =   1 ' b 0 ;     w r _ c y c l e [       3 9 ]   =   1 ' b 1 ;     a d d r _ r o m [       3 9 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       3 9 ] = ' h 0 0 0 0 0 0 3 d ;  
         r d _ c y c l e [       4 0 ]   =   1 ' b 1 ;     w r _ c y c l e [       4 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       4 0 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [       4 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       4 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       4 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       4 1 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [       4 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       4 2 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 2 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 2 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [       4 2 ] = ' h 0 0 0 0 0 0 1 7 ;  
         r d _ c y c l e [       4 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       4 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       4 3 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       4 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       4 4 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 4 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 4 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       4 4 ] = ' h 0 0 0 0 0 0 0 2 ;  
         r d _ c y c l e [       4 5 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 5 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 5 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       4 5 ] = ' h 0 0 0 0 0 0 2 5 ;  
         r d _ c y c l e [       4 6 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 6 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 6 ] = ' h 0 0 0 0 0 0 3 0 ;     w r _ d a t a _ r o m [       4 6 ] = ' h 0 0 0 0 0 0 0 1 ;  
         r d _ c y c l e [       4 7 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 7 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 7 ] = ' h 0 0 0 0 0 0 0 4 ;     w r _ d a t a _ r o m [       4 7 ] = ' h 0 0 0 0 0 0 0 6 ;  
         r d _ c y c l e [       4 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 8 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 8 ] = ' h 0 0 0 0 0 0 2 0 ;     w r _ d a t a _ r o m [       4 8 ] = ' h 0 0 0 0 0 0 0 d ;  
         r d _ c y c l e [       4 9 ]   =   1 ' b 0 ;     w r _ c y c l e [       4 9 ]   =   1 ' b 1 ;     a d d r _ r o m [       4 9 ] = ' h 0 0 0 0 0 0 2 4 ;     w r _ d a t a _ r o m [       4 9 ] = ' h 0 0 0 0 0 0 1 7 ;  
         r d _ c y c l e [       5 0 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 0 ] = ' h 0 0 0 0 0 0 3 c ;     w r _ d a t a _ r o m [       5 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 1 ]   =   1 ' b 0 ;     w r _ c y c l e [       5 1 ]   =   1 ' b 1 ;     a d d r _ r o m [       5 1 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       5 1 ] = ' h 0 0 0 0 0 0 2 9 ;  
         r d _ c y c l e [       5 2 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 2 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 2 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       5 2 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 3 ] = ' h 0 0 0 0 0 0 1 4 ;     w r _ d a t a _ r o m [       5 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 4 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 4 ] = ' h 0 0 0 0 0 0 0 8 ;     w r _ d a t a _ r o m [       5 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 5 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 5 ] = ' h 0 0 0 0 0 0 3 4 ;     w r _ d a t a _ r o m [       5 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 6 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 6 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 6 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       5 6 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       5 7 ]   =   1 ' b 0 ;     w r _ c y c l e [       5 7 ]   =   1 ' b 1 ;     a d d r _ r o m [       5 7 ] = ' h 0 0 0 0 0 0 2 0 ;     w r _ d a t a _ r o m [       5 7 ] = ' h 0 0 0 0 0 0 0 9 ;  
         r d _ c y c l e [       5 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       5 8 ]   =   1 ' b 1 ;     a d d r _ r o m [       5 8 ] = ' h 0 0 0 0 0 0 0 8 ;     w r _ d a t a _ r o m [       5 8 ] = ' h 0 0 0 0 0 0 1 0 ;  
         r d _ c y c l e [       5 9 ]   =   1 ' b 1 ;     w r _ c y c l e [       5 9 ]   =   1 ' b 0 ;     a d d r _ r o m [       5 9 ] = ' h 0 0 0 0 0 0 2 8 ;     w r _ d a t a _ r o m [       5 9 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 0 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 0 ]   =   1 ' b 1 ;     a d d r _ r o m [       6 0 ] = ' h 0 0 0 0 0 0 2 4 ;     w r _ d a t a _ r o m [       6 0 ] = ' h 0 0 0 0 0 0 0 b ;  
         r d _ c y c l e [       6 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       6 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 1 ] = ' h 0 0 0 0 0 0 3 c ;     w r _ d a t a _ r o m [       6 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 2 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 2 ]   =   1 ' b 1 ;     a d d r _ r o m [       6 2 ] = ' h 0 0 0 0 0 0 3 0 ;     w r _ d a t a _ r o m [       6 2 ] = ' h 0 0 0 0 0 0 0 4 ;  
         r d _ c y c l e [       6 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       6 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 3 ] = ' h 0 0 0 0 0 0 2 c ;     w r _ d a t a _ r o m [       6 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         / /   1 6   s i l e n c e   c y c l e s  
         r d _ c y c l e [       6 4 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 4 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 5 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 5 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 6 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 6 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 6 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 6 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 7 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 7 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 8 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 8 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 8 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       6 9 ]   =   1 ' b 0 ;     w r _ c y c l e [       6 9 ]   =   1 ' b 0 ;     a d d r _ r o m [       6 9 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       6 9 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 0 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 0 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 1 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 1 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 2 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 2 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 2 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 2 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 3 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 3 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 4 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 4 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 5 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 5 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 6 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 6 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 6 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 6 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 7 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 7 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 8 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 8 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 8 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 8 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       7 9 ]   =   1 ' b 0 ;     w r _ c y c l e [       7 9 ]   =   1 ' b 0 ;     a d d r _ r o m [       7 9 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       7 9 ] = ' h 0 0 0 0 0 0 0 0 ;  
         / /   1 6   s e q u e n c e   r e a d   c y c l e s  
         r d _ c y c l e [       8 0 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 0 ] = ' h 0 0 0 0 0 0 0 0 ;     w r _ d a t a _ r o m [       8 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 1 ] = ' h 0 0 0 0 0 0 0 4 ;     w r _ d a t a _ r o m [       8 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 2 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 2 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 2 ] = ' h 0 0 0 0 0 0 0 8 ;     w r _ d a t a _ r o m [       8 2 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 3 ] = ' h 0 0 0 0 0 0 0 c ;     w r _ d a t a _ r o m [       8 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 4 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 4 ] = ' h 0 0 0 0 0 0 1 0 ;     w r _ d a t a _ r o m [       8 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 5 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 5 ] = ' h 0 0 0 0 0 0 1 4 ;     w r _ d a t a _ r o m [       8 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 6 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 6 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 6 ] = ' h 0 0 0 0 0 0 1 8 ;     w r _ d a t a _ r o m [       8 6 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 7 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 7 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 7 ] = ' h 0 0 0 0 0 0 1 c ;     w r _ d a t a _ r o m [       8 7 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 8 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 8 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 8 ] = ' h 0 0 0 0 0 0 2 0 ;     w r _ d a t a _ r o m [       8 8 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       8 9 ]   =   1 ' b 1 ;     w r _ c y c l e [       8 9 ]   =   1 ' b 0 ;     a d d r _ r o m [       8 9 ] = ' h 0 0 0 0 0 0 2 4 ;     w r _ d a t a _ r o m [       8 9 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 0 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 0 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 0 ] = ' h 0 0 0 0 0 0 2 8 ;     w r _ d a t a _ r o m [       9 0 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 1 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 1 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 1 ] = ' h 0 0 0 0 0 0 2 c ;     w r _ d a t a _ r o m [       9 1 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 2 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 2 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 2 ] = ' h 0 0 0 0 0 0 3 0 ;     w r _ d a t a _ r o m [       9 2 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 3 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 3 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 3 ] = ' h 0 0 0 0 0 0 3 4 ;     w r _ d a t a _ r o m [       9 3 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 4 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 4 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 4 ] = ' h 0 0 0 0 0 0 3 8 ;     w r _ d a t a _ r o m [       9 4 ] = ' h 0 0 0 0 0 0 0 0 ;  
         r d _ c y c l e [       9 5 ]   =   1 ' b 1 ;     w r _ c y c l e [       9 5 ]   =   1 ' b 0 ;     a d d r _ r o m [       9 5 ] = ' h 0 0 0 0 0 0 3 c ;     w r _ d a t a _ r o m [       9 5 ] = ' h 0 0 0 0 0 0 0 0 ;  
 e n d  
  
 i n i t i a l   b e g i n  
         v a l i d a t i o n _ d a t a [         0 ]   =   ' h 0 0 0 0 0 0 2 9 ;    
         v a l i d a t i o n _ d a t a [         1 ]   =   ' h 0 0 0 0 0 0 0 6 ;    
         v a l i d a t i o n _ d a t a [         2 ]   =   ' h 0 0 0 0 0 0 1 0 ;    
         v a l i d a t i o n _ d a t a [         3 ]   =   ' h 0 0 0 0 0 0 1 2 ;    
         v a l i d a t i o n _ d a t a [         4 ]   =   ' h 0 0 0 0 0 0 0 e ;    
         v a l i d a t i o n _ d a t a [         5 ]   =   ' h 0 0 0 0 0 0 0 4 ;    
         v a l i d a t i o n _ d a t a [         6 ]   =   ' h 0 0 0 0 0 0 1 0 ;    
         v a l i d a t i o n _ d a t a [         7 ]   =   ' h 0 0 0 0 0 0 1 7 ;    
         v a l i d a t i o n _ d a t a [         8 ]   =   ' h 0 0 0 0 0 0 0 9 ;    
         v a l i d a t i o n _ d a t a [         9 ]   =   ' h 0 0 0 0 0 0 0 b ;    
         v a l i d a t i o n _ d a t a [       1 0 ]   =   ' h 0 0 0 0 0 0 1 e ;    
         v a l i d a t i o n _ d a t a [       1 1 ]   =   ' h 0 0 0 0 0 0 2 6 ;    
         v a l i d a t i o n _ d a t a [       1 2 ]   =   ' h 0 0 0 0 0 0 0 4 ;    
         v a l i d a t i o n _ d a t a [       1 3 ]   =   ' h 0 0 0 0 0 0 3 e ;    
         v a l i d a t i o n _ d a t a [       1 4 ]   =   ' h 0 0 0 0 0 0 0 2 ;    
         v a l i d a t i o n _ d a t a [       1 5 ]   =   ' h 0 0 0 0 0 0 1 4 ;    
  
 e n d  
  
  
 r e g   c l k   =   1 ' b 1 ,   r s t   =   1 ' b 1 ;  
 i n i t i a l   # 4   r s t   =   1 ' b 0 ;  
 a l w a y s     # 1   c l k   =   ~ c l k ;  
  
 w i r e     m i s s ;  
 w i r e   [ 3 1 : 0 ]   r d _ d a t a ;  
 r e g     [ 3 1 : 0 ]   i n d e x   =   0 ,   w r _ d a t a   =   0 ,   a d d r   =   0 ;  
 r e g     r d _ r e q   =   1 ' b 0 ,   w r _ r e q   =   1 ' b 0 ;  
 r e g   r d _ r e q _ f f   =   1 ' b 0 ,   m i s s _ f f   =   1 ' b 0 ;  
 r e g   [ 3 1 : 0 ]   v a l i d a t i o n _ c o u n t   =   0 ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )   b e g i n  
                 r d _ r e q _ f f   < =   1 ' b 0 ;  
                 m i s s _ f f       < =   1 ' b 0 ;  
         e n d   e l s e   b e g i n  
                 r d _ r e q _ f f   < =   r d _ r e q ;  
                 m i s s _ f f       < =   m i s s ;  
         e n d  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )   b e g i n  
                 v a l i d a t i o n _ c o u n t   < =   0 ;  
         e n d   e l s e   b e g i n  
                 i f ( v a l i d a t i o n _ c o u n t > = ` D A T A _ C O U N T )   b e g i n  
                         v a l i d a t i o n _ c o u n t   < =   ' h f f f f f f f f ;  
                 e n d   e l s e   i f ( r d _ r e q _ f f   & &   ( i n d e x > ( 4 * ` D A T A _ C O U N T ) ) )   b e g i n  
                         i f ( ~ m i s s _ f f )   b e g i n  
                                 i f ( v a l i d a t i o n _ d a t a [ v a l i d a t i o n _ c o u n t ] = = r d _ d a t a )  
                                         v a l i d a t i o n _ c o u n t   < =   v a l i d a t i o n _ c o u n t + 1 ;  
                                 e l s e  
                                         v a l i d a t i o n _ c o u n t   < =   0 ;  
                         e n d  
                 e n d   e l s e   b e g i n  
                         v a l i d a t i o n _ c o u n t   < =   0 ;  
                 e n d  
         e n d  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )   b e g i n  
                 i n d e x       < =   0 ;  
                 w r _ d a t a   < =   0 ;  
                 a d d r         < =   0 ;  
                 r d _ r e q     < =   1 ' b 0 ;  
                 w r _ r e q     < =   1 ' b 0 ;  
         e n d   e l s e   b e g i n  
                 i f ( ~ m i s s )   b e g i n  
                         i f ( i n d e x < ` R D W R _ C O U N T )   b e g i n  
                                 i f ( w r _ c y c l e [ i n d e x ] )   b e g i n  
                                         r d _ r e q     < =   1 ' b 0 ;  
                                         w r _ r e q     < =   1 ' b 1 ;  
                                 e n d   e l s e   i f ( r d _ c y c l e [ i n d e x ] )   b e g i n  
                                         w r _ d a t a   < =   0 ;  
                                         r d _ r e q     < =   1 ' b 1 ;  
                                         w r _ r e q     < =   1 ' b 0 ;  
                                 e n d   e l s e   b e g i n  
                                         w r _ d a t a   < =   0 ;  
                                         r d _ r e q     < =   1 ' b 0 ;  
                                         w r _ r e q     < =   1 ' b 0 ;  
                                 e n d  
                                 w r _ d a t a   < =   w r _ d a t a _ r o m [ i n d e x ] ;  
                                 a d d r         < =   a d d r _ r o m [ i n d e x ] ;  
                                 i n d e x   < =   i n d e x   +   1 ;  
                         e n d   e l s e   b e g i n  
                                 w r _ d a t a   < =   0 ;  
                                 a d d r         < =   0 ;  
                                 r d _ r e q     < =   1 ' b 0 ;  
                                 w r _ r e q     < =   1 ' b 0 ;  
                         e n d  
                 e n d  
         e n d  
  
 c a c h e   # (  
         . L I N E _ A D D R _ L E N     (   3                           ) ,  
         . S E T _ A D D R _ L E N       (   2                           ) ,  
         . T A G _ A D D R _ L E N       (   1 2                         ) ,  
         . W A Y _ C N T                 (   3                           )  
 )   c a c h e _ t e s t _ i n s t a n c e   (  
         . c l k                         (   c l k                       ) ,  
         . r s t                         (   r s t                       ) ,  
         . m i s s                       (   m i s s                     ) ,  
         . a d d r                       (   a d d r                     ) ,  
         . r d _ r e q                   (   r d _ r e q                 ) ,  
         . r d _ d a t a                 (   r d _ d a t a               ) ,  
         . w r _ r e q                   (   w r _ r e q                 ) ,  
         . w r _ d a t a                 (   w r _ d a t a               )  
 ) ;  
  
 e n d m o d u l e  
  
 