�� 
 m o d u l e   m e m   # (                                       / /    
         p a r a m e t e r     A D D R _ L E N     =   1 1       / /    
 )   (  
         i n p u t     c l k ,   r s t ,  
         i n p u t     [ A D D R _ L E N - 1 : 0 ]   a d d r ,   / /   m e m o r y   a d d r e s s  
         o u t p u t   r e g   [ 3 1 : 0 ]   r d _ d a t a ,     / /   d a t a   r e a d   o u t  
         i n p u t     w r _ r e q ,  
         i n p u t     [ 3 1 : 0 ]   w r _ d a t a               / /   d a t a   w r i t e   i n  
 ) ;  
 l o c a l p a r a m   M E M _ S I Z E   =   1 < < A D D R _ L E N ;  
 r e g   [ 3 1 : 0 ]   r a m _ c e l l   [ M E M _ S I Z E ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k   o r   p o s e d g e   r s t )  
         i f ( r s t )  
                 r d _ d a t a   < =   0 ;  
         e l s e  
                 r d _ d a t a   < =   r a m _ c e l l [ a d d r ] ;  
  
 a l w a y s   @   ( p o s e d g e   c l k )  
         i f ( w r _ r e q )    
                 r a m _ c e l l [ a d d r ]   < =   w r _ d a t a ;  
  
 i n i t i a l   b e g i n  
         / /   d s t   m a t r i x   C  
         r a m _ c e l l [               0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 9 1 f c d 2 e ;  
         r a m _ c e l l [               1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e f f 3 d 5 2 0 ;  
         r a m _ c e l l [               2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b d 8 4 7 b 8 4 ;  
         r a m _ c e l l [               3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 0 e 9 c 8 4 b ;  
         r a m _ c e l l [               4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 8 5 7 0 3 2 0 ;  
         r a m _ c e l l [               5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b b 7 6 e 8 4 1 ;  
         r a m _ c e l l [               6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 4 f 2 6 2 9 ;  
         r a m _ c e l l [               7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 e b f 2 1 7 0 ;  
         r a m _ c e l l [               8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 b 5 f 3 d b ;  
         r a m _ c e l l [               9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 e e 5 7 1 5 6 ;  
         r a m _ c e l l [             1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 c 8 b e 7 f ;  
         r a m _ c e l l [             1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 b a 0 7 f 2 0 ;  
         r a m _ c e l l [             1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 d 6 7 3 9 3 d ;  
         r a m _ c e l l [             1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 d 7 e 7 3 5 ;  
         r a m _ c e l l [             1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 a a f 7 b 7 ;  
         r a m _ c e l l [             1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 8 6 7 3 7 1 7 ;  
         r a m _ c e l l [             1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 9 c 9 1 a 8 4 ;  
         r a m _ c e l l [             1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 b a 2 6 2 4 3 ;  
         r a m _ c e l l [             1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 9 5 9 f 6 3 8 ;  
         r a m _ c e l l [             1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d b 6 3 2 4 9 5 ;  
         r a m _ c e l l [             2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 9 e b c c d 5 ;  
         r a m _ c e l l [             2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 0 2 a f 6 7 b ;  
         r a m _ c e l l [             2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f 5 2 f 3 0 0 ;  
         r a m _ c e l l [             2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 0 c e 2 b 2 a ;  
         r a m _ c e l l [             2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 d 5 0 1 e 8 d ;  
         r a m _ c e l l [             2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 c 3 6 d 6 e 9 ;  
         r a m _ c e l l [             2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 6 5 e 7 5 0 2 ;  
         r a m _ c e l l [             2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 0 b 8 a 7 b d ;  
         r a m _ c e l l [             2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b c 5 4 0 a d 7 ;  
         r a m _ c e l l [             2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 8 9 4 8 9 9 d ;  
         r a m _ c e l l [             3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f b 0 6 7 4 5 7 ;  
         r a m _ c e l l [             3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d f 1 7 e 9 2 4 ;  
         r a m _ c e l l [             3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 1 9 b 4 1 1 f ;  
         r a m _ c e l l [             3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c f d d 3 8 f a ;  
         r a m _ c e l l [             3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c d e 0 5 e 8 2 ;  
         r a m _ c e l l [             3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 4 b 1 6 6 3 8 ;  
         r a m _ c e l l [             3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 4 4 7 d 1 1 2 ;  
         r a m _ c e l l [             3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 4 7 6 0 b 2 4 ;  
         r a m _ c e l l [             3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 9 f c f 8 b e ;  
         r a m _ c e l l [             3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 b 4 3 4 2 8 2 ;  
         r a m _ c e l l [             4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 0 8 f c 7 8 5 ;  
         r a m _ c e l l [             4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 1 d 5 c c e d ;  
         r a m _ c e l l [             4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 0 4 1 6 5 5 d ;  
         r a m _ c e l l [             4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 5 a b 9 0 d 0 ;  
         r a m _ c e l l [             4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 7 b 6 1 c d a ;  
         r a m _ c e l l [             4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 3 1 9 5 1 4 1 ;  
         r a m _ c e l l [             4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 3 5 b a 4 5 f ;  
         r a m _ c e l l [             4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a f 8 c 5 4 2 c ;  
         r a m _ c e l l [             4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 9 d 6 9 8 1 a ;  
         r a m _ c e l l [             4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 3 a 3 3 c 1 1 ;  
         r a m _ c e l l [             5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 b 0 0 3 2 2 7 ;  
         r a m _ c e l l [             5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 7 8 d 1 2 1 ;  
         r a m _ c e l l [             5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 e 7 c e 8 7 d ;  
         r a m _ c e l l [             5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 4 b c 2 f d 2 ;  
         r a m _ c e l l [             5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 8 e 1 8 0 f 3 ;  
         r a m _ c e l l [             5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 d 5 c 9 1 5 1 ;  
         r a m _ c e l l [             5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 0 e f 5 5 c f ;  
         r a m _ c e l l [             5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 2 8 e 8 d b 9 ;  
         r a m _ c e l l [             5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f 5 5 e 2 3 f ;  
         r a m _ c e l l [             5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 7 e 3 9 c c 4 ;  
         r a m _ c e l l [             6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 c c f 1 4 5 c ;  
         r a m _ c e l l [             6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d e d 4 7 3 b 6 ;  
         r a m _ c e l l [             6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 b 9 c e 2 f 9 ;  
         r a m _ c e l l [             6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f c 8 a 4 e 3 e ;  
         r a m _ c e l l [             6 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 e e 6 0 a 4 b ;  
         r a m _ c e l l [             6 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 f 3 5 d 8 d ;  
         r a m _ c e l l [             6 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 b 1 1 5 7 e 7 ;  
         r a m _ c e l l [             6 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 9 e b 2 4 6 6 ;  
         r a m _ c e l l [             6 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f e e 7 c 7 3 f ;  
         r a m _ c e l l [             6 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 4 c 4 e 9 9 3 ;  
         r a m _ c e l l [             7 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 4 4 c b 1 5 f ;  
         r a m _ c e l l [             7 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 3 d 3 1 9 9 0 ;  
         r a m _ c e l l [             7 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 f f b d d a b ;  
         r a m _ c e l l [             7 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 2 4 5 e 3 9 3 ;  
         r a m _ c e l l [             7 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 9 0 d 5 e b 7 ;  
         r a m _ c e l l [             7 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a a 9 5 1 c 6 2 ;  
         r a m _ c e l l [             7 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 9 f 1 3 d f 5 ;  
         r a m _ c e l l [             7 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d b c 3 b 5 0 a ;  
         r a m _ c e l l [             7 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 2 8 a d f 7 6 ;  
         r a m _ c e l l [             7 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c b 4 3 7 a 6 1 ;  
         r a m _ c e l l [             8 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 9 5 3 8 7 6 7 ;  
         r a m _ c e l l [             8 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 b 8 0 7 9 6 5 ;  
         r a m _ c e l l [             8 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 7 9 9 6 6 e e ;  
         r a m _ c e l l [             8 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 3 9 a 1 8 9 7 ;  
         r a m _ c e l l [             8 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 f a e 9 9 2 2 ;  
         r a m _ c e l l [             8 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 e 2 8 a c d b ;  
         r a m _ c e l l [             8 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 c d 5 0 4 3 d ;  
         r a m _ c e l l [             8 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 b 9 0 4 f e 5 ;  
         r a m _ c e l l [             8 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 e 0 2 c 1 0 d ;  
         r a m _ c e l l [             8 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 5 0 6 b 8 7 9 ;  
         r a m _ c e l l [             9 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 2 c 9 0 5 8 5 ;  
         r a m _ c e l l [             9 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 3 c 7 a 1 f d ;  
         r a m _ c e l l [             9 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d b 0 9 8 9 5 a ;  
         r a m _ c e l l [             9 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 1 a c 5 1 9 b ;  
         r a m _ c e l l [             9 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 5 1 e d 5 d 1 ;  
         r a m _ c e l l [             9 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 6 8 1 3 e 5 ;  
         r a m _ c e l l [             9 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a f b 8 a a 7 1 ;  
         r a m _ c e l l [             9 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 f 5 c 6 9 c 9 ;  
         r a m _ c e l l [             9 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 0 9 3 1 4 c ;  
         r a m _ c e l l [             9 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 e 7 9 5 9 b b ;  
         r a m _ c e l l [           1 0 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 2 d 5 9 e 4 ;  
         r a m _ c e l l [           1 0 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 f e a f 8 3 a ;  
         r a m _ c e l l [           1 0 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 f 2 0 7 8 0 0 ;  
         r a m _ c e l l [           1 0 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c f 3 0 4 8 c 0 ;  
         r a m _ c e l l [           1 0 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 9 3 8 8 a f 6 ;  
         r a m _ c e l l [           1 0 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 4 4 1 5 0 8 6 ;  
         r a m _ c e l l [           1 0 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c d 2 4 f 5 d 5 ;  
         r a m _ c e l l [           1 0 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 1 c b e a a 6 ;  
         r a m _ c e l l [           1 0 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 0 9 2 2 5 3 9 ;  
         r a m _ c e l l [           1 0 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 9 d 4 4 e 7 b ;  
         r a m _ c e l l [           1 1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 5 5 c f 4 a 9 ;  
         r a m _ c e l l [           1 1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 d 6 c 7 6 7 5 ;  
         r a m _ c e l l [           1 1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 7 c b 6 3 1 2 ;  
         r a m _ c e l l [           1 1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 d 8 f 4 1 2 9 ;  
         r a m _ c e l l [           1 1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 8 0 b e 9 2 1 ;  
         r a m _ c e l l [           1 1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e f 6 b 5 2 c 4 ;  
         r a m _ c e l l [           1 1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 0 9 8 7 c a 9 ;  
         r a m _ c e l l [           1 1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 2 6 2 5 9 8 0 ;  
         r a m _ c e l l [           1 1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 2 c 1 f 7 c 6 ;  
         r a m _ c e l l [           1 1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 5 e 2 a 4 d 5 ;  
         r a m _ c e l l [           1 2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e c 5 2 8 3 e c ;  
         r a m _ c e l l [           1 2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 4 6 a 1 1 0 8 ;  
         r a m _ c e l l [           1 2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 4 8 a b 1 9 6 ;  
         r a m _ c e l l [           1 2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 c 2 b 6 7 f f ;  
         r a m _ c e l l [           1 2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 3 7 7 3 8 9 f ;  
         r a m _ c e l l [           1 2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 4 8 8 b b 0 e ;  
         r a m _ c e l l [           1 2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 b 7 6 3 c b 3 ;  
         r a m _ c e l l [           1 2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 2 d f 7 9 3 2 ;  
         r a m _ c e l l [           1 2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f d 7 0 2 5 1 1 ;  
         r a m _ c e l l [           1 2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 2 5 e 1 a 4 c ;  
         r a m _ c e l l [           1 3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 5 3 6 2 1 f 7 ;  
         r a m _ c e l l [           1 3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 1 d 0 d b 2 ;  
         r a m _ c e l l [           1 3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 f b 9 7 2 1 2 ;  
         r a m _ c e l l [           1 3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 9 2 d 1 2 0 b ;  
         r a m _ c e l l [           1 3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 0 f 7 2 6 9 5 ;  
         r a m _ c e l l [           1 3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 a 7 a 7 a 5 6 ;  
         r a m _ c e l l [           1 3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 f e 7 d 3 d e ;  
         r a m _ c e l l [           1 3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 3 c c e a c 0 ;  
         r a m _ c e l l [           1 3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 e 7 c 1 1 5 9 ;  
         r a m _ c e l l [           1 3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 1 1 e f 3 2 7 ;  
         r a m _ c e l l [           1 4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 8 7 d 3 0 d e ;  
         r a m _ c e l l [           1 4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 d 2 c 0 1 8 8 ;  
         r a m _ c e l l [           1 4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 0 6 2 d 4 5 3 ;  
         r a m _ c e l l [           1 4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 3 2 c b b 0 d ;  
         r a m _ c e l l [           1 4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 9 0 7 7 1 8 f ;  
         r a m _ c e l l [           1 4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 0 b b 9 2 f 7 ;  
         r a m _ c e l l [           1 4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 f 8 a f 5 3 2 ;  
         r a m _ c e l l [           1 4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b f 2 2 2 f a f ;  
         r a m _ c e l l [           1 4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 1 9 7 0 7 2 3 ;  
         r a m _ c e l l [           1 4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 4 f 2 5 d 9 e ;  
         r a m _ c e l l [           1 5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 3 0 c a 2 5 b ;  
         r a m _ c e l l [           1 5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 1 b 3 d f b 7 ;  
         r a m _ c e l l [           1 5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 5 d 2 3 1 c b ;  
         r a m _ c e l l [           1 5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 7 2 a 5 0 b 1 ;  
         r a m _ c e l l [           1 5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 b 1 7 0 8 b 4 ;  
         r a m _ c e l l [           1 5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 9 0 b 8 1 3 f ;  
         r a m _ c e l l [           1 5 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 1 d d 2 2 5 1 ;  
         r a m _ c e l l [           1 5 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 4 b 4 2 c 9 7 ;  
         r a m _ c e l l [           1 5 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f d e d 9 c 7 f ;  
         r a m _ c e l l [           1 5 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 6 1 b a 6 a b ;  
         r a m _ c e l l [           1 6 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e f 8 0 6 f e c ;  
         r a m _ c e l l [           1 6 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 a d a 2 9 3 c ;  
         r a m _ c e l l [           1 6 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 b 7 d 5 0 b d ;  
         r a m _ c e l l [           1 6 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c d 8 3 c 2 4 c ;  
         r a m _ c e l l [           1 6 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c a 1 4 f 2 b e ;  
         r a m _ c e l l [           1 6 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 6 d f d b a e ;  
         r a m _ c e l l [           1 6 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 1 3 b 3 b 4 8 ;  
         r a m _ c e l l [           1 6 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d d 4 3 f 8 f f ;  
         r a m _ c e l l [           1 6 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 8 5 d 9 9 e 3 ;  
         r a m _ c e l l [           1 6 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 9 6 8 d e 0 9 ;  
         r a m _ c e l l [           1 7 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 8 a 5 4 5 5 f ;  
         r a m _ c e l l [           1 7 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 0 5 0 1 4 b 7 ;  
         r a m _ c e l l [           1 7 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 3 d f 9 e 3 c ;  
         r a m _ c e l l [           1 7 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 7 9 7 a 6 e b ;  
         r a m _ c e l l [           1 7 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 4 a f b 8 d 0 ;  
         r a m _ c e l l [           1 7 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 f b c c a c d ;  
         r a m _ c e l l [           1 7 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 8 2 b 9 d 4 6 ;  
         r a m _ c e l l [           1 7 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 5 9 c c 1 5 9 ;  
         r a m _ c e l l [           1 7 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 b 4 c b a 8 6 ;  
         r a m _ c e l l [           1 7 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 8 6 d f a 8 6 ;  
         r a m _ c e l l [           1 8 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 c 2 9 e 2 f e ;  
         r a m _ c e l l [           1 8 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 6 b 1 0 b b 5 ;  
         r a m _ c e l l [           1 8 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f 1 2 b 2 f 0 ;  
         r a m _ c e l l [           1 8 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 c 4 5 f 5 e 3 ;  
         r a m _ c e l l [           1 8 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 7 b d 4 4 1 b ;  
         r a m _ c e l l [           1 8 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 2 8 d f 2 e 4 ;  
         r a m _ c e l l [           1 8 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f e 0 6 c c 4 2 ;  
         r a m _ c e l l [           1 8 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 6 e 6 1 9 4 4 ;  
         r a m _ c e l l [           1 8 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 c 8 b f 2 7 f ;  
         r a m _ c e l l [           1 8 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 c 3 f 2 5 4 c ;  
         r a m _ c e l l [           1 9 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 3 a 0 7 6 c 0 ;  
         r a m _ c e l l [           1 9 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 4 a 3 2 8 6 7 ;  
         r a m _ c e l l [           1 9 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 c 1 2 5 6 c c ;  
         r a m _ c e l l [           1 9 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 8 c 2 3 6 5 5 ;  
         r a m _ c e l l [           1 9 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 0 5 4 2 7 1 6 ;  
         r a m _ c e l l [           1 9 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 5 a 7 f 5 b d ;  
         r a m _ c e l l [           1 9 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 1 c 3 7 b 9 9 ;  
         r a m _ c e l l [           1 9 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 2 1 1 0 5 7 3 ;  
         r a m _ c e l l [           1 9 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a 2 2 7 6 c 4 b ;  
         r a m _ c e l l [           1 9 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 3 4 2 4 1 3 2 ;  
         r a m _ c e l l [           2 0 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 3 b e d 9 0 9 ;  
         r a m _ c e l l [           2 0 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 5 4 b 8 3 a 8 ;  
         r a m _ c e l l [           2 0 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 3 2 b c e 7 9 ;  
         r a m _ c e l l [           2 0 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 f e 3 2 7 6 9 ;  
         r a m _ c e l l [           2 0 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 2 8 9 c b 2 4 ;  
         r a m _ c e l l [           2 0 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a c 9 8 d 5 7 8 ;  
         r a m _ c e l l [           2 0 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 1 f 6 6 1 e 1 ;  
         r a m _ c e l l [           2 0 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 4 f c 7 9 d 2 ;  
         r a m _ c e l l [           2 0 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 c 0 b c 6 2 1 ;  
         r a m _ c e l l [           2 0 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 6 b 7 7 7 4 0 0 ;  
         r a m _ c e l l [           2 1 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 5 5 1 9 2 1 e ;  
         r a m _ c e l l [           2 1 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 c 5 1 0 a 8 f ;  
         r a m _ c e l l [           2 1 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a b e 3 7 f 1 8 ;  
         r a m _ c e l l [           2 1 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h a e 4 3 9 c 3 7 ;  
         r a m _ c e l l [           2 1 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 1 4 6 f d a 5 ;  
         r a m _ c e l l [           2 1 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b d e a e 0 5 4 ;  
         r a m _ c e l l [           2 1 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 8 a d 8 3 b 7 ;  
         r a m _ c e l l [           2 1 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 8 4 e f f 7 5 ;  
         r a m _ c e l l [           2 1 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 4 1 c 1 7 2 9 ;  
         r a m _ c e l l [           2 1 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 0 5 1 a 7 4 7 ;  
         r a m _ c e l l [           2 2 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 3 2 9 8 0 1 7 ;  
         r a m _ c e l l [           2 2 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e a f 9 a 6 e 0 ;  
         r a m _ c e l l [           2 2 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 8 5 f a 6 2 1 ;  
         r a m _ c e l l [           2 2 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 b 7 b a 8 f 5 ;  
         r a m _ c e l l [           2 2 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 d 5 a 1 b 7 1 ;  
         r a m _ c e l l [           2 2 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 5 c d 2 d d f ;  
         r a m _ c e l l [           2 2 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 d a 8 2 0 a f ;  
         r a m _ c e l l [           2 2 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 d 2 7 d a e e ;  
         r a m _ c e l l [           2 2 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 5 1 b 1 0 b d ;  
         r a m _ c e l l [           2 2 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 5 d 7 5 7 2 5 ;  
         r a m _ c e l l [           2 3 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 9 1 e c a 7 f ;  
         r a m _ c e l l [           2 3 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 8 8 0 b 3 9 c ;  
         r a m _ c e l l [           2 3 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 7 8 2 f b 0 4 d ;  
         r a m _ c e l l [           2 3 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 3 8 c f 6 5 f ;  
         r a m _ c e l l [           2 3 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 1 f c 7 5 6 0 ;  
         r a m _ c e l l [           2 3 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h d 7 2 9 7 9 f 0 ;  
         r a m _ c e l l [           2 3 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h c 5 e 0 5 1 0 d ;  
         r a m _ c e l l [           2 3 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 6 9 7 1 b e e ;  
         r a m _ c e l l [           2 3 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e b 1 7 3 9 0 f ;  
         r a m _ c e l l [           2 3 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 9 8 0 a d f 5 b ;  
         r a m _ c e l l [           2 4 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 a c d f b 6 f ;  
         r a m _ c e l l [           2 4 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 3 6 3 8 0 8 b ;  
         r a m _ c e l l [           2 4 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 1 7 f 4 7 7 d ;  
         r a m _ c e l l [           2 4 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 9 5 3 4 4 1 b ;  
         r a m _ c e l l [           2 4 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f 4 9 0 b 0 6 d ;  
         r a m _ c e l l [           2 4 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 5 8 b 8 5 a 4 3 ;  
         r a m _ c e l l [           2 4 6 ]   =   3 2 ' h 0 ;     / /   3 2 ' h f b f 0 9 b b 5 ;  
         r a m _ c e l l [           2 4 7 ]   =   3 2 ' h 0 ;     / /   3 2 ' h e 9 8 f 5 9 2 e ;  
         r a m _ c e l l [           2 4 8 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 4 8 f 8 7 d a a ;  
         r a m _ c e l l [           2 4 9 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 1 b 9 c b b 7 a ;  
         r a m _ c e l l [           2 5 0 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 7 4 3 6 1 0 2 ;  
         r a m _ c e l l [           2 5 1 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 0 0 8 e 7 c 5 5 ;  
         r a m _ c e l l [           2 5 2 ]   =   3 2 ' h 0 ;     / /   3 2 ' h b 1 f 4 f 2 7 0 ;  
         r a m _ c e l l [           2 5 3 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 8 f 8 9 6 a c 8 ;  
         r a m _ c e l l [           2 5 4 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 3 5 3 e 3 8 5 5 ;  
         r a m _ c e l l [           2 5 5 ]   =   3 2 ' h 0 ;     / /   3 2 ' h 2 a 6 0 d 3 4 4 ;  
         / /   s r c   m a t r i x   A  
         r a m _ c e l l [           2 5 6 ]   =   3 2 ' h 5 8 2 b 6 9 f 0 ;  
         r a m _ c e l l [           2 5 7 ]   =   3 2 ' h 5 1 c e 9 6 8 9 ;  
         r a m _ c e l l [           2 5 8 ]   =   3 2 ' h 6 d f 6 0 a 3 0 ;  
         r a m _ c e l l [           2 5 9 ]   =   3 2 ' h 3 1 a a f 4 f 8 ;  
         r a m _ c e l l [           2 6 0 ]   =   3 2 ' h a 3 4 7 b a 1 5 ;  
         r a m _ c e l l [           2 6 1 ]   =   3 2 ' h 6 d d d e a e 0 ;  
         r a m _ c e l l [           2 6 2 ]   =   3 2 ' h d 3 9 c 4 6 1 0 ;  
         r a m _ c e l l [           2 6 3 ]   =   3 2 ' h 8 3 7 1 3 e 5 9 ;  
         r a m _ c e l l [           2 6 4 ]   =   3 2 ' h 9 3 f e 2 7 5 d ;  
         r a m _ c e l l [           2 6 5 ]   =   3 2 ' h 9 e 1 0 5 2 7 3 ;  
         r a m _ c e l l [           2 6 6 ]   =   3 2 ' h 5 9 6 5 2 9 e 2 ;  
         r a m _ c e l l [           2 6 7 ]   =   3 2 ' h 5 9 4 c 2 6 6 d ;  
         r a m _ c e l l [           2 6 8 ]   =   3 2 ' h a 4 3 9 6 7 1 e ;  
         r a m _ c e l l [           2 6 9 ]   =   3 2 ' h f 4 c 7 b c b 8 ;  
         r a m _ c e l l [           2 7 0 ]   =   3 2 ' h d b d 7 c 5 5 e ;  
         r a m _ c e l l [           2 7 1 ]   =   3 2 ' h 8 4 7 3 4 d 5 5 ;  
         r a m _ c e l l [           2 7 2 ]   =   3 2 ' h 1 9 e 0 6 2 4 0 ;  
         r a m _ c e l l [           2 7 3 ]   =   3 2 ' h 5 0 c c 0 4 3 8 ;  
         r a m _ c e l l [           2 7 4 ]   =   3 2 ' h b c c 7 2 4 b 0 ;  
         r a m _ c e l l [           2 7 5 ]   =   3 2 ' h 2 d b b e a 6 a ;  
         r a m _ c e l l [           2 7 6 ]   =   3 2 ' h d b 1 2 4 9 8 a ;  
         r a m _ c e l l [           2 7 7 ]   =   3 2 ' h a e a a e 8 6 1 ;  
         r a m _ c e l l [           2 7 8 ]   =   3 2 ' h 8 f d 3 4 0 a 8 ;  
         r a m _ c e l l [           2 7 9 ]   =   3 2 ' h c 5 c a c f e 0 ;  
         r a m _ c e l l [           2 8 0 ]   =   3 2 ' h 0 3 7 9 2 e 3 2 ;  
         r a m _ c e l l [           2 8 1 ]   =   3 2 ' h e 6 a 0 7 6 b a ;  
         r a m _ c e l l [           2 8 2 ]   =   3 2 ' h 9 f 3 e 0 2 e 5 ;  
         r a m _ c e l l [           2 8 3 ]   =   3 2 ' h 9 f 0 4 c b e f ;  
         r a m _ c e l l [           2 8 4 ]   =   3 2 ' h b 6 e 1 0 f d b ;  
         r a m _ c e l l [           2 8 5 ]   =   3 2 ' h c 9 7 1 e 0 2 9 ;  
         r a m _ c e l l [           2 8 6 ]   =   3 2 ' h f 8 5 e 4 3 5 e ;  
         r a m _ c e l l [           2 8 7 ]   =   3 2 ' h 6 1 b e 4 5 6 a ;  
         r a m _ c e l l [           2 8 8 ]   =   3 2 ' h 0 1 6 4 4 4 9 2 ;  
         r a m _ c e l l [           2 8 9 ]   =   3 2 ' h 4 0 0 0 a 1 7 2 ;  
         r a m _ c e l l [           2 9 0 ]   =   3 2 ' h c 8 6 a 9 2 c 8 ;  
         r a m _ c e l l [           2 9 1 ]   =   3 2 ' h b 8 0 b f 8 1 5 ;  
         r a m _ c e l l [           2 9 2 ]   =   3 2 ' h 1 e 9 6 2 7 8 7 ;  
         r a m _ c e l l [           2 9 3 ]   =   3 2 ' h 3 5 2 f 9 f 8 a ;  
         r a m _ c e l l [           2 9 4 ]   =   3 2 ' h 8 6 0 6 3 a 2 6 ;  
         r a m _ c e l l [           2 9 5 ]   =   3 2 ' h 3 4 1 6 2 1 6 6 ;  
         r a m _ c e l l [           2 9 6 ]   =   3 2 ' h 9 2 5 0 a 5 e a ;  
         r a m _ c e l l [           2 9 7 ]   =   3 2 ' h 2 7 e 7 8 0 f 2 ;  
         r a m _ c e l l [           2 9 8 ]   =   3 2 ' h c d 0 4 8 d 2 a ;  
         r a m _ c e l l [           2 9 9 ]   =   3 2 ' h 6 2 6 c d 2 b 4 ;  
         r a m _ c e l l [           3 0 0 ]   =   3 2 ' h 2 8 4 e b 6 d d ;  
         r a m _ c e l l [           3 0 1 ]   =   3 2 ' h 5 0 e 4 c 5 f 4 ;  
         r a m _ c e l l [           3 0 2 ]   =   3 2 ' h 5 0 8 9 a b 1 6 ;  
         r a m _ c e l l [           3 0 3 ]   =   3 2 ' h c 1 e 9 2 8 7 8 ;  
         r a m _ c e l l [           3 0 4 ]   =   3 2 ' h 2 6 c 9 c a 0 0 ;  
         r a m _ c e l l [           3 0 5 ]   =   3 2 ' h 8 8 1 0 b b 4 9 ;  
         r a m _ c e l l [           3 0 6 ]   =   3 2 ' h e e 6 a 9 1 c b ;  
         r a m _ c e l l [           3 0 7 ]   =   3 2 ' h 0 3 1 5 9 b 2 3 ;  
         r a m _ c e l l [           3 0 8 ]   =   3 2 ' h 0 6 d f 1 4 a 7 ;  
         r a m _ c e l l [           3 0 9 ]   =   3 2 ' h f 5 3 a 8 9 d 3 ;  
         r a m _ c e l l [           3 1 0 ]   =   3 2 ' h 0 c 7 9 f a 6 8 ;  
         r a m _ c e l l [           3 1 1 ]   =   3 2 ' h 7 2 7 e d 4 8 b ;  
         r a m _ c e l l [           3 1 2 ]   =   3 2 ' h 7 c c 0 5 a 9 7 ;  
         r a m _ c e l l [           3 1 3 ]   =   3 2 ' h f a 8 c 2 d b d ;  
         r a m _ c e l l [           3 1 4 ]   =   3 2 ' h 4 f 3 6 7 5 8 e ;  
         r a m _ c e l l [           3 1 5 ]   =   3 2 ' h d 7 b 8 1 a 7 d ;  
         r a m _ c e l l [           3 1 6 ]   =   3 2 ' h d 8 9 d b d 6 9 ;  
         r a m _ c e l l [           3 1 7 ]   =   3 2 ' h 3 f f a 3 9 b 8 ;  
         r a m _ c e l l [           3 1 8 ]   =   3 2 ' h d 2 d b 4 5 8 f ;  
         r a m _ c e l l [           3 1 9 ]   =   3 2 ' h 9 4 9 3 9 a 0 3 ;  
         r a m _ c e l l [           3 2 0 ]   =   3 2 ' h d 5 3 7 8 6 e 2 ;  
         r a m _ c e l l [           3 2 1 ]   =   3 2 ' h e 4 f a f f f c ;  
         r a m _ c e l l [           3 2 2 ]   =   3 2 ' h 5 8 1 c b 2 b 9 ;  
         r a m _ c e l l [           3 2 3 ]   =   3 2 ' h f 8 4 d 6 4 5 5 ;  
         r a m _ c e l l [           3 2 4 ]   =   3 2 ' h b 8 a d d 6 e 4 ;  
         r a m _ c e l l [           3 2 5 ]   =   3 2 ' h 1 7 4 7 6 5 4 1 ;  
         r a m _ c e l l [           3 2 6 ]   =   3 2 ' h e 9 4 d 5 2 c f ;  
         r a m _ c e l l [           3 2 7 ]   =   3 2 ' h 6 0 e 0 5 d d c ;  
         r a m _ c e l l [           3 2 8 ]   =   3 2 ' h 6 f 3 9 1 e 6 6 ;  
         r a m _ c e l l [           3 2 9 ]   =   3 2 ' h 3 e 9 d 9 b 0 f ;  
         r a m _ c e l l [           3 3 0 ]   =   3 2 ' h 3 2 f e 0 9 a 5 ;  
         r a m _ c e l l [           3 3 1 ]   =   3 2 ' h 9 d e 7 3 9 c 7 ;  
         r a m _ c e l l [           3 3 2 ]   =   3 2 ' h b 3 1 f 1 4 6 7 ;  
         r a m _ c e l l [           3 3 3 ]   =   3 2 ' h 1 b 5 6 4 c 5 9 ;  
         r a m _ c e l l [           3 3 4 ]   =   3 2 ' h d 4 e 5 8 1 e c ;  
         r a m _ c e l l [           3 3 5 ]   =   3 2 ' h 2 5 8 4 a f e 6 ;  
         r a m _ c e l l [           3 3 6 ]   =   3 2 ' h e 5 f 6 c 4 1 c ;  
         r a m _ c e l l [           3 3 7 ]   =   3 2 ' h c a f 8 e c 0 9 ;  
         r a m _ c e l l [           3 3 8 ]   =   3 2 ' h 4 c 2 7 b 1 2 7 ;  
         r a m _ c e l l [           3 3 9 ]   =   3 2 ' h 7 e 5 7 e 6 0 a ;  
         r a m _ c e l l [           3 4 0 ]   =   3 2 ' h 1 5 2 1 3 7 1 b ;  
         r a m _ c e l l [           3 4 1 ]   =   3 2 ' h c 5 8 1 b 7 1 3 ;  
         r a m _ c e l l [           3 4 2 ]   =   3 2 ' h 5 7 5 4 9 5 7 d ;  
         r a m _ c e l l [           3 4 3 ]   =   3 2 ' h e 7 c 9 e 0 8 b ;  
         r a m _ c e l l [           3 4 4 ]   =   3 2 ' h 7 8 9 3 a e 4 7 ;  
         r a m _ c e l l [           3 4 5 ]   =   3 2 ' h 3 f a 3 1 4 a 3 ;  
         r a m _ c e l l [           3 4 6 ]   =   3 2 ' h e a 7 2 6 f d 3 ;  
         r a m _ c e l l [           3 4 7 ]   =   3 2 ' h 0 f 9 8 1 1 6 1 ;  
         r a m _ c e l l [           3 4 8 ]   =   3 2 ' h e 8 2 b f 8 b 3 ;  
         r a m _ c e l l [           3 4 9 ]   =   3 2 ' h e b 4 4 9 9 0 f ;  
         r a m _ c e l l [           3 5 0 ]   =   3 2 ' h c 6 3 6 9 0 2 f ;  
         r a m _ c e l l [           3 5 1 ]   =   3 2 ' h 6 6 3 6 e b 7 3 ;  
         r a m _ c e l l [           3 5 2 ]   =   3 2 ' h a f a 3 2 5 6 a ;  
         r a m _ c e l l [           3 5 3 ]   =   3 2 ' h 6 9 6 b 2 4 7 9 ;  
         r a m _ c e l l [           3 5 4 ]   =   3 2 ' h b f 9 b f a 5 e ;  
         r a m _ c e l l [           3 5 5 ]   =   3 2 ' h 3 4 1 1 f 2 e 5 ;  
         r a m _ c e l l [           3 5 6 ]   =   3 2 ' h 8 f 9 2 4 7 b 3 ;  
         r a m _ c e l l [           3 5 7 ]   =   3 2 ' h 6 c 6 c 1 f 2 4 ;  
         r a m _ c e l l [           3 5 8 ]   =   3 2 ' h 5 7 9 4 a 1 d 2 ;  
         r a m _ c e l l [           3 5 9 ]   =   3 2 ' h b 4 d 9 7 a 5 2 ;  
         r a m _ c e l l [           3 6 0 ]   =   3 2 ' h e f d 0 2 7 6 7 ;  
         r a m _ c e l l [           3 6 1 ]   =   3 2 ' h 0 a 0 f 8 8 4 1 ;  
         r a m _ c e l l [           3 6 2 ]   =   3 2 ' h 0 3 3 d 1 4 7 6 ;  
         r a m _ c e l l [           3 6 3 ]   =   3 2 ' h 3 5 4 c 6 8 1 6 ;  
         r a m _ c e l l [           3 6 4 ]   =   3 2 ' h 6 7 9 b 7 1 b 7 ;  
         r a m _ c e l l [           3 6 5 ]   =   3 2 ' h a b 3 1 3 8 1 9 ;  
         r a m _ c e l l [           3 6 6 ]   =   3 2 ' h 7 f 0 5 7 f 1 8 ;  
         r a m _ c e l l [           3 6 7 ]   =   3 2 ' h 6 8 b b c 5 1 4 ;  
         r a m _ c e l l [           3 6 8 ]   =   3 2 ' h 2 d b 2 0 6 3 c ;  
         r a m _ c e l l [           3 6 9 ]   =   3 2 ' h 9 f f 1 f c e 0 ;  
         r a m _ c e l l [           3 7 0 ]   =   3 2 ' h e 7 a 4 8 5 0 9 ;  
         r a m _ c e l l [           3 7 1 ]   =   3 2 ' h b 0 8 6 d 7 9 5 ;  
         r a m _ c e l l [           3 7 2 ]   =   3 2 ' h 5 9 5 7 5 a 3 7 ;  
         r a m _ c e l l [           3 7 3 ]   =   3 2 ' h 7 4 a 2 9 9 d 6 ;  
         r a m _ c e l l [           3 7 4 ]   =   3 2 ' h 8 8 a c b a b 4 ;  
         r a m _ c e l l [           3 7 5 ]   =   3 2 ' h a 2 c 5 2 f a 7 ;  
         r a m _ c e l l [           3 7 6 ]   =   3 2 ' h 4 b 5 a d 5 a a ;  
         r a m _ c e l l [           3 7 7 ]   =   3 2 ' h 6 2 7 1 5 9 9 d ;  
         r a m _ c e l l [           3 7 8 ]   =   3 2 ' h a d 9 c e 3 b 3 ;  
         r a m _ c e l l [           3 7 9 ]   =   3 2 ' h a 7 4 2 a f f 1 ;  
         r a m _ c e l l [           3 8 0 ]   =   3 2 ' h b f 6 6 c 9 3 a ;  
         r a m _ c e l l [           3 8 1 ]   =   3 2 ' h 0 6 d c 4 0 3 a ;  
         r a m _ c e l l [           3 8 2 ]   =   3 2 ' h 7 a 8 4 8 3 7 b ;  
         r a m _ c e l l [           3 8 3 ]   =   3 2 ' h 0 d c b a d 0 1 ;  
         r a m _ c e l l [           3 8 4 ]   =   3 2 ' h d f e b f d e 6 ;  
         r a m _ c e l l [           3 8 5 ]   =   3 2 ' h 3 7 b 5 c a b d ;  
         r a m _ c e l l [           3 8 6 ]   =   3 2 ' h 1 6 3 8 1 1 2 d ;  
         r a m _ c e l l [           3 8 7 ]   =   3 2 ' h 9 2 c 8 7 d e 9 ;  
         r a m _ c e l l [           3 8 8 ]   =   3 2 ' h 2 a 9 4 7 5 e c ;  
         r a m _ c e l l [           3 8 9 ]   =   3 2 ' h b d d a e 7 b 4 ;  
         r a m _ c e l l [           3 9 0 ]   =   3 2 ' h 9 d d 4 b 5 8 0 ;  
         r a m _ c e l l [           3 9 1 ]   =   3 2 ' h 0 9 c b 5 1 b c ;  
         r a m _ c e l l [           3 9 2 ]   =   3 2 ' h f 5 1 0 5 c 9 4 ;  
         r a m _ c e l l [           3 9 3 ]   =   3 2 ' h 9 9 d e 9 d 0 4 ;  
         r a m _ c e l l [           3 9 4 ]   =   3 2 ' h 7 7 1 8 c b e a ;  
         r a m _ c e l l [           3 9 5 ]   =   3 2 ' h 0 0 d 1 7 5 8 7 ;  
         r a m _ c e l l [           3 9 6 ]   =   3 2 ' h e 0 7 9 e 8 4 8 ;  
         r a m _ c e l l [           3 9 7 ]   =   3 2 ' h 9 f b 0 4 5 3 e ;  
         r a m _ c e l l [           3 9 8 ]   =   3 2 ' h c 2 7 9 6 1 b e ;  
         r a m _ c e l l [           3 9 9 ]   =   3 2 ' h 5 2 7 4 9 5 9 a ;  
         r a m _ c e l l [           4 0 0 ]   =   3 2 ' h b 0 f 9 c 5 0 7 ;  
         r a m _ c e l l [           4 0 1 ]   =   3 2 ' h 0 8 9 f 5 1 3 a ;  
         r a m _ c e l l [           4 0 2 ]   =   3 2 ' h 9 a c c f 5 d 0 ;  
         r a m _ c e l l [           4 0 3 ]   =   3 2 ' h 1 f f 6 8 c c 3 ;  
         r a m _ c e l l [           4 0 4 ]   =   3 2 ' h 7 d 9 2 9 6 4 e ;  
         r a m _ c e l l [           4 0 5 ]   =   3 2 ' h 3 e d e 9 b 9 1 ;  
         r a m _ c e l l [           4 0 6 ]   =   3 2 ' h 6 7 a 7 5 e 6 e ;  
         r a m _ c e l l [           4 0 7 ]   =   3 2 ' h f 5 9 1 4 b 1 d ;  
         r a m _ c e l l [           4 0 8 ]   =   3 2 ' h 8 a d 9 5 2 7 d ;  
         r a m _ c e l l [           4 0 9 ]   =   3 2 ' h d 6 d 8 8 8 c 2 ;  
         r a m _ c e l l [           4 1 0 ]   =   3 2 ' h 9 b 2 8 a e f b ;  
         r a m _ c e l l [           4 1 1 ]   =   3 2 ' h 2 0 d 7 f a 0 2 ;  
         r a m _ c e l l [           4 1 2 ]   =   3 2 ' h a 9 0 9 9 8 9 a ;  
         r a m _ c e l l [           4 1 3 ]   =   3 2 ' h e b e 5 3 b b b ;  
         r a m _ c e l l [           4 1 4 ]   =   3 2 ' h 7 f f 4 e 8 8 0 ;  
         r a m _ c e l l [           4 1 5 ]   =   3 2 ' h 2 6 0 e e e b 4 ;  
         r a m _ c e l l [           4 1 6 ]   =   3 2 ' h 5 4 2 5 0 7 1 6 ;  
         r a m _ c e l l [           4 1 7 ]   =   3 2 ' h 3 8 0 7 4 c 3 3 ;  
         r a m _ c e l l [           4 1 8 ]   =   3 2 ' h b 4 d 0 9 c 1 8 ;  
         r a m _ c e l l [           4 1 9 ]   =   3 2 ' h c d a 6 2 4 7 f ;  
         r a m _ c e l l [           4 2 0 ]   =   3 2 ' h 7 2 5 4 8 b 1 9 ;  
         r a m _ c e l l [           4 2 1 ]   =   3 2 ' h b 5 1 d 6 a d 6 ;  
         r a m _ c e l l [           4 2 2 ]   =   3 2 ' h 2 0 f 6 1 0 4 a ;  
         r a m _ c e l l [           4 2 3 ]   =   3 2 ' h 6 4 8 c c 9 b 9 ;  
         r a m _ c e l l [           4 2 4 ]   =   3 2 ' h 9 6 4 8 6 8 9 f ;  
         r a m _ c e l l [           4 2 5 ]   =   3 2 ' h 0 9 0 c 7 c 7 8 ;  
         r a m _ c e l l [           4 2 6 ]   =   3 2 ' h 4 f 6 d a e 9 d ;  
         r a m _ c e l l [           4 2 7 ]   =   3 2 ' h 2 6 7 e 1 2 5 a ;  
         r a m _ c e l l [           4 2 8 ]   =   3 2 ' h f 6 7 f 7 4 1 8 ;  
         r a m _ c e l l [           4 2 9 ]   =   3 2 ' h c 8 3 7 1 8 c 8 ;  
         r a m _ c e l l [           4 3 0 ]   =   3 2 ' h 5 9 3 1 f 2 9 6 ;  
         r a m _ c e l l [           4 3 1 ]   =   3 2 ' h 8 4 4 5 0 b 4 c ;  
         r a m _ c e l l [           4 3 2 ]   =   3 2 ' h 5 1 6 c 2 0 7 6 ;  
         r a m _ c e l l [           4 3 3 ]   =   3 2 ' h 8 e 4 3 8 3 3 8 ;  
         r a m _ c e l l [           4 3 4 ]   =   3 2 ' h e 7 a 9 b 7 d b ;  
         r a m _ c e l l [           4 3 5 ]   =   3 2 ' h 8 c 6 1 1 d 8 9 ;  
         r a m _ c e l l [           4 3 6 ]   =   3 2 ' h d 9 c 8 e 0 b 2 ;  
         r a m _ c e l l [           4 3 7 ]   =   3 2 ' h 6 5 f 7 c a 7 4 ;  
         r a m _ c e l l [           4 3 8 ]   =   3 2 ' h 6 2 0 0 1 3 2 9 ;  
         r a m _ c e l l [           4 3 9 ]   =   3 2 ' h 1 b 0 9 3 1 6 8 ;  
         r a m _ c e l l [           4 4 0 ]   =   3 2 ' h 0 d e 5 6 4 e 4 ;  
         r a m _ c e l l [           4 4 1 ]   =   3 2 ' h 8 4 8 6 5 3 8 1 ;  
         r a m _ c e l l [           4 4 2 ]   =   3 2 ' h f 5 9 9 d 6 1 8 ;  
         r a m _ c e l l [           4 4 3 ]   =   3 2 ' h 6 f 6 f a 5 4 a ;  
         r a m _ c e l l [           4 4 4 ]   =   3 2 ' h 3 a b 3 7 4 c 6 ;  
         r a m _ c e l l [           4 4 5 ]   =   3 2 ' h 7 e 7 2 0 5 0 d ;  
         r a m _ c e l l [           4 4 6 ]   =   3 2 ' h 4 6 9 b f 8 a a ;  
         r a m _ c e l l [           4 4 7 ]   =   3 2 ' h 0 1 5 b 6 a e a ;  
         r a m _ c e l l [           4 4 8 ]   =   3 2 ' h b d 9 4 e 8 7 3 ;  
         r a m _ c e l l [           4 4 9 ]   =   3 2 ' h 7 c 2 0 c 9 8 c ;  
         r a m _ c e l l [           4 5 0 ]   =   3 2 ' h 9 7 0 6 f 1 0 9 ;  
         r a m _ c e l l [           4 5 1 ]   =   3 2 ' h 2 3 3 2 1 4 b 1 ;  
         r a m _ c e l l [           4 5 2 ]   =   3 2 ' h 8 4 6 d 2 e 2 a ;  
         r a m _ c e l l [           4 5 3 ]   =   3 2 ' h 7 0 3 c 5 5 1 f ;  
         r a m _ c e l l [           4 5 4 ]   =   3 2 ' h 2 5 3 b 1 d a d ;  
         r a m _ c e l l [           4 5 5 ]   =   3 2 ' h 6 7 e a 6 2 c 1 ;  
         r a m _ c e l l [           4 5 6 ]   =   3 2 ' h 3 1 9 2 7 4 3 1 ;  
         r a m _ c e l l [           4 5 7 ]   =   3 2 ' h b 6 f f 9 a 1 4 ;  
         r a m _ c e l l [           4 5 8 ]   =   3 2 ' h f 8 1 e 2 c 7 c ;  
         r a m _ c e l l [           4 5 9 ]   =   3 2 ' h a 6 7 d 7 3 3 9 ;  
         r a m _ c e l l [           4 6 0 ]   =   3 2 ' h 7 7 6 8 d 0 7 8 ;  
         r a m _ c e l l [           4 6 1 ]   =   3 2 ' h 5 2 8 9 e c e d ;  
         r a m _ c e l l [           4 6 2 ]   =   3 2 ' h 8 f 7 c 1 6 d 8 ;  
         r a m _ c e l l [           4 6 3 ]   =   3 2 ' h 1 8 9 6 0 f b f ;  
         r a m _ c e l l [           4 6 4 ]   =   3 2 ' h e 1 4 0 e e 3 4 ;  
         r a m _ c e l l [           4 6 5 ]   =   3 2 ' h d 5 6 2 5 8 9 f ;  
         r a m _ c e l l [           4 6 6 ]   =   3 2 ' h 7 4 d 4 2 0 9 0 ;  
         r a m _ c e l l [           4 6 7 ]   =   3 2 ' h a 2 7 d a 2 0 5 ;  
         r a m _ c e l l [           4 6 8 ]   =   3 2 ' h 2 2 3 2 7 b b a ;  
         r a m _ c e l l [           4 6 9 ]   =   3 2 ' h 2 6 c c c 2 2 f ;  
         r a m _ c e l l [           4 7 0 ]   =   3 2 ' h c 8 c c 9 9 9 7 ;  
         r a m _ c e l l [           4 7 1 ]   =   3 2 ' h 9 3 8 b d b 0 e ;  
         r a m _ c e l l [           4 7 2 ]   =   3 2 ' h 5 b 0 8 c 9 0 c ;  
         r a m _ c e l l [           4 7 3 ]   =   3 2 ' h 6 d a 9 e 2 6 0 ;  
         r a m _ c e l l [           4 7 4 ]   =   3 2 ' h 7 e 9 0 d 0 9 4 ;  
         r a m _ c e l l [           4 7 5 ]   =   3 2 ' h 7 0 a d e 8 b 0 ;  
         r a m _ c e l l [           4 7 6 ]   =   3 2 ' h 0 9 2 1 0 2 0 7 ;  
         r a m _ c e l l [           4 7 7 ]   =   3 2 ' h 9 d f a b b 5 c ;  
         r a m _ c e l l [           4 7 8 ]   =   3 2 ' h c b b e a a f 7 ;  
         r a m _ c e l l [           4 7 9 ]   =   3 2 ' h 2 4 8 5 5 b 4 e ;  
         r a m _ c e l l [           4 8 0 ]   =   3 2 ' h d 8 a f c b 1 a ;  
         r a m _ c e l l [           4 8 1 ]   =   3 2 ' h 4 7 9 2 f 8 f 3 ;  
         r a m _ c e l l [           4 8 2 ]   =   3 2 ' h b 0 1 9 3 4 5 9 ;  
         r a m _ c e l l [           4 8 3 ]   =   3 2 ' h a 8 5 b b 2 a 7 ;  
         r a m _ c e l l [           4 8 4 ]   =   3 2 ' h e 0 9 e a 0 f 7 ;  
         r a m _ c e l l [           4 8 5 ]   =   3 2 ' h 9 0 d 1 7 d 0 6 ;  
         r a m _ c e l l [           4 8 6 ]   =   3 2 ' h a f c 8 f 2 d e ;  
         r a m _ c e l l [           4 8 7 ]   =   3 2 ' h 9 d f 2 d 4 e 8 ;  
         r a m _ c e l l [           4 8 8 ]   =   3 2 ' h 5 6 8 5 a 8 1 6 ;  
         r a m _ c e l l [           4 8 9 ]   =   3 2 ' h 4 2 b a 1 4 f c ;  
         r a m _ c e l l [           4 9 0 ]   =   3 2 ' h 6 2 0 2 b 3 7 d ;  
         r a m _ c e l l [           4 9 1 ]   =   3 2 ' h 5 a b 3 8 d e 1 ;  
         r a m _ c e l l [           4 9 2 ]   =   3 2 ' h d 4 e b e 4 6 e ;  
         r a m _ c e l l [           4 9 3 ]   =   3 2 ' h f f d b a 9 6 7 ;  
         r a m _ c e l l [           4 9 4 ]   =   3 2 ' h 6 7 2 b 7 8 1 c ;  
         r a m _ c e l l [           4 9 5 ]   =   3 2 ' h a e 0 3 d 0 0 8 ;  
         r a m _ c e l l [           4 9 6 ]   =   3 2 ' h 0 8 5 c d 7 7 8 ;  
         r a m _ c e l l [           4 9 7 ]   =   3 2 ' h 5 1 d 8 7 4 7 6 ;  
         r a m _ c e l l [           4 9 8 ]   =   3 2 ' h f 9 b 3 f 0 8 c ;  
         r a m _ c e l l [           4 9 9 ]   =   3 2 ' h b d 7 d c b f b ;  
         r a m _ c e l l [           5 0 0 ]   =   3 2 ' h 6 c c 3 2 2 0 3 ;  
         r a m _ c e l l [           5 0 1 ]   =   3 2 ' h 2 7 a e 0 d d 1 ;  
         r a m _ c e l l [           5 0 2 ]   =   3 2 ' h f 8 2 0 7 d 7 7 ;  
         r a m _ c e l l [           5 0 3 ]   =   3 2 ' h 8 f f 3 6 f 1 3 ;  
         r a m _ c e l l [           5 0 4 ]   =   3 2 ' h c 4 e 9 3 c 8 f ;  
         r a m _ c e l l [           5 0 5 ]   =   3 2 ' h f f 8 b 6 7 6 9 ;  
         r a m _ c e l l [           5 0 6 ]   =   3 2 ' h 4 d 5 3 6 5 1 3 ;  
         r a m _ c e l l [           5 0 7 ]   =   3 2 ' h d d 9 8 4 e 3 8 ;  
         r a m _ c e l l [           5 0 8 ]   =   3 2 ' h 7 f 6 2 c a e d ;  
         r a m _ c e l l [           5 0 9 ]   =   3 2 ' h 7 3 3 d 9 a 2 a ;  
         r a m _ c e l l [           5 1 0 ]   =   3 2 ' h 1 8 3 1 8 a 1 0 ;  
         r a m _ c e l l [           5 1 1 ]   =   3 2 ' h 1 6 c 8 b 2 c 6 ;  
         / /   s r c   m a t r i x   B  
         r a m _ c e l l [           5 1 2 ]   =   3 2 ' h 7 d 0 f 8 3 f 4 ;  
         r a m _ c e l l [           5 1 3 ]   =   3 2 ' h b e c 2 e b 7 0 ;  
         r a m _ c e l l [           5 1 4 ]   =   3 2 ' h c 6 7 e 3 4 b 2 ;  
         r a m _ c e l l [           5 1 5 ]   =   3 2 ' h 9 b f 6 a 1 a 9 ;  
         r a m _ c e l l [           5 1 6 ]   =   3 2 ' h 3 3 d f 3 6 9 e ;  
         r a m _ c e l l [           5 1 7 ]   =   3 2 ' h 3 5 b c 7 8 3 a ;  
         r a m _ c e l l [           5 1 8 ]   =   3 2 ' h b c 8 d e b 4 c ;  
         r a m _ c e l l [           5 1 9 ]   =   3 2 ' h 2 0 9 d b 1 5 1 ;  
         r a m _ c e l l [           5 2 0 ]   =   3 2 ' h c c 3 f 8 1 9 9 ;  
         r a m _ c e l l [           5 2 1 ]   =   3 2 ' h d 0 3 d 6 5 3 9 ;  
         r a m _ c e l l [           5 2 2 ]   =   3 2 ' h c a 4 e 6 6 1 f ;  
         r a m _ c e l l [           5 2 3 ]   =   3 2 ' h 6 3 e 0 6 f d 1 ;  
         r a m _ c e l l [           5 2 4 ]   =   3 2 ' h f 2 1 e 9 2 1 9 ;  
         r a m _ c e l l [           5 2 5 ]   =   3 2 ' h 3 2 0 f a 9 1 d ;  
         r a m _ c e l l [           5 2 6 ]   =   3 2 ' h 4 1 9 d e 3 7 b ;  
         r a m _ c e l l [           5 2 7 ]   =   3 2 ' h 1 0 2 9 4 c 9 b ;  
         r a m _ c e l l [           5 2 8 ]   =   3 2 ' h 1 1 8 5 1 4 a 2 ;  
         r a m _ c e l l [           5 2 9 ]   =   3 2 ' h 5 7 4 8 d 1 3 8 ;  
         r a m _ c e l l [           5 3 0 ]   =   3 2 ' h 6 1 f 1 1 4 7 4 ;  
         r a m _ c e l l [           5 3 1 ]   =   3 2 ' h 3 5 b b b b 0 e ;  
         r a m _ c e l l [           5 3 2 ]   =   3 2 ' h 1 6 9 7 1 e 0 2 ;  
         r a m _ c e l l [           5 3 3 ]   =   3 2 ' h d 3 6 9 a 6 b 0 ;  
         r a m _ c e l l [           5 3 4 ]   =   3 2 ' h 8 2 3 b e d 9 9 ;  
         r a m _ c e l l [           5 3 5 ]   =   3 2 ' h 0 9 b 2 b a 3 d ;  
         r a m _ c e l l [           5 3 6 ]   =   3 2 ' h 0 9 4 6 0 f b 1 ;  
         r a m _ c e l l [           5 3 7 ]   =   3 2 ' h 6 3 e c d 2 5 c ;  
         r a m _ c e l l [           5 3 8 ]   =   3 2 ' h d 2 c 8 a c 1 8 ;  
         r a m _ c e l l [           5 3 9 ]   =   3 2 ' h 9 4 5 c 8 7 f 6 ;  
         r a m _ c e l l [           5 4 0 ]   =   3 2 ' h 1 c 0 d e 2 2 e ;  
         r a m _ c e l l [           5 4 1 ]   =   3 2 ' h f 5 4 a f b d 1 ;  
         r a m _ c e l l [           5 4 2 ]   =   3 2 ' h 9 c 2 2 3 d f 4 ;  
         r a m _ c e l l [           5 4 3 ]   =   3 2 ' h 9 c 5 e 3 0 e b ;  
         r a m _ c e l l [           5 4 4 ]   =   3 2 ' h 0 a b 0 8 9 e 1 ;  
         r a m _ c e l l [           5 4 5 ]   =   3 2 ' h 9 7 5 7 e c 5 3 ;  
         r a m _ c e l l [           5 4 6 ]   =   3 2 ' h 3 2 f 0 f 6 c f ;  
         r a m _ c e l l [           5 4 7 ]   =   3 2 ' h f e c f a a 7 1 ;  
         r a m _ c e l l [           5 4 8 ]   =   3 2 ' h 5 7 8 8 9 0 7 2 ;  
         r a m _ c e l l [           5 4 9 ]   =   3 2 ' h 1 6 9 a c 0 3 4 ;  
         r a m _ c e l l [           5 5 0 ]   =   3 2 ' h 5 d 3 c d f c e ;  
         r a m _ c e l l [           5 5 1 ]   =   3 2 ' h e c a e d 1 7 7 ;  
         r a m _ c e l l [           5 5 2 ]   =   3 2 ' h 0 a 7 6 2 3 c 8 ;  
         r a m _ c e l l [           5 5 3 ]   =   3 2 ' h d 4 2 d 9 3 5 5 ;  
         r a m _ c e l l [           5 5 4 ]   =   3 2 ' h 8 6 a e e 6 b 4 ;  
         r a m _ c e l l [           5 5 5 ]   =   3 2 ' h e f 4 0 3 b 9 3 ;  
         r a m _ c e l l [           5 5 6 ]   =   3 2 ' h 6 4 c 7 a 1 a f ;  
         r a m _ c e l l [           5 5 7 ]   =   3 2 ' h e 4 e 4 4 7 9 3 ;  
         r a m _ c e l l [           5 5 8 ]   =   3 2 ' h 2 c a 8 8 4 e 4 ;  
         r a m _ c e l l [           5 5 9 ]   =   3 2 ' h 8 4 a b a b 8 d ;  
         r a m _ c e l l [           5 6 0 ]   =   3 2 ' h 0 d 8 3 7 f 3 e ;  
         r a m _ c e l l [           5 6 1 ]   =   3 2 ' h 6 a b 1 f 0 f 6 ;  
         r a m _ c e l l [           5 6 2 ]   =   3 2 ' h 1 a 0 e 5 4 7 9 ;  
         r a m _ c e l l [           5 6 3 ]   =   3 2 ' h 8 f f 6 4 a e 3 ;  
         r a m _ c e l l [           5 6 4 ]   =   3 2 ' h 4 7 a 9 e 8 8 e ;  
         r a m _ c e l l [           5 6 5 ]   =   3 2 ' h e 4 1 a 0 1 f e ;  
         r a m _ c e l l [           5 6 6 ]   =   3 2 ' h 0 7 1 1 1 3 f f ;  
         r a m _ c e l l [           5 6 7 ]   =   3 2 ' h d d e 5 5 a 7 4 ;  
         r a m _ c e l l [           5 6 8 ]   =   3 2 ' h f 2 2 f e 5 1 2 ;  
         r a m _ c e l l [           5 6 9 ]   =   3 2 ' h 5 3 6 5 a 9 e d ;  
         r a m _ c e l l [           5 7 0 ]   =   3 2 ' h 6 a d 6 7 a 6 8 ;  
         r a m _ c e l l [           5 7 1 ]   =   3 2 ' h 2 d 8 9 5 8 c 8 ;  
         r a m _ c e l l [           5 7 2 ]   =   3 2 ' h b 4 7 4 d 3 f 4 ;  
         r a m _ c e l l [           5 7 3 ]   =   3 2 ' h f 9 5 2 1 b e d ;  
         r a m _ c e l l [           5 7 4 ]   =   3 2 ' h d a 3 3 b c 1 7 ;  
         r a m _ c e l l [           5 7 5 ]   =   3 2 ' h e e e 3 2 9 4 8 ;  
         r a m _ c e l l [           5 7 6 ]   =   3 2 ' h 8 f 3 4 f 2 b f ;  
         r a m _ c e l l [           5 7 7 ]   =   3 2 ' h b 6 5 1 5 8 5 7 ;  
         r a m _ c e l l [           5 7 8 ]   =   3 2 ' h a 5 a b f e f e ;  
         r a m _ c e l l [           5 7 9 ]   =   3 2 ' h c 8 9 f e c 0 3 ;  
         r a m _ c e l l [           5 8 0 ]   =   3 2 ' h 5 0 5 0 9 0 e 3 ;  
         r a m _ c e l l [           5 8 1 ]   =   3 2 ' h 6 d 8 6 9 c 0 d ;  
         r a m _ c e l l [           5 8 2 ]   =   3 2 ' h 7 9 4 1 5 e 3 3 ;  
         r a m _ c e l l [           5 8 3 ]   =   3 2 ' h d 0 9 1 3 a 8 3 ;  
         r a m _ c e l l [           5 8 4 ]   =   3 2 ' h 3 c 1 8 8 d 0 f ;  
         r a m _ c e l l [           5 8 5 ]   =   3 2 ' h 7 e 8 a d 9 b 5 ;  
         r a m _ c e l l [           5 8 6 ]   =   3 2 ' h a 8 9 0 5 6 7 a ;  
         r a m _ c e l l [           5 8 7 ]   =   3 2 ' h c 9 f c d b a 8 ;  
         r a m _ c e l l [           5 8 8 ]   =   3 2 ' h d 7 4 7 3 1 2 6 ;  
         r a m _ c e l l [           5 8 9 ]   =   3 2 ' h 5 6 3 c a 0 1 7 ;  
         r a m _ c e l l [           5 9 0 ]   =   3 2 ' h d 5 f a d 3 b 4 ;  
         r a m _ c e l l [           5 9 1 ]   =   3 2 ' h 5 3 1 5 0 8 6 b ;  
         r a m _ c e l l [           5 9 2 ]   =   3 2 ' h 1 4 5 c 7 7 1 1 ;  
         r a m _ c e l l [           5 9 3 ]   =   3 2 ' h 6 7 5 e a 8 9 1 ;  
         r a m _ c e l l [           5 9 4 ]   =   3 2 ' h e 7 d b 0 6 7 0 ;  
         r a m _ c e l l [           5 9 5 ]   =   3 2 ' h 7 5 d 2 b 1 b a ;  
         r a m _ c e l l [           5 9 6 ]   =   3 2 ' h 5 e d e 6 9 6 c ;  
         r a m _ c e l l [           5 9 7 ]   =   3 2 ' h e 9 1 1 c 2 e 8 ;  
         r a m _ c e l l [           5 9 8 ]   =   3 2 ' h 1 6 5 0 0 7 6 2 ;  
         r a m _ c e l l [           5 9 9 ]   =   3 2 ' h e 8 a 5 0 7 0 8 ;  
         r a m _ c e l l [           6 0 0 ]   =   3 2 ' h 1 0 c 1 9 4 9 2 ;  
         r a m _ c e l l [           6 0 1 ]   =   3 2 ' h 3 8 b 9 7 4 e 4 ;  
         r a m _ c e l l [           6 0 2 ]   =   3 2 ' h 7 4 c 7 f 7 b 9 ;  
         r a m _ c e l l [           6 0 3 ]   =   3 2 ' h 3 d 3 7 1 b 0 6 ;  
         r a m _ c e l l [           6 0 4 ]   =   3 2 ' h 7 3 c 5 9 c d 9 ;  
         r a m _ c e l l [           6 0 5 ]   =   3 2 ' h c 2 f 5 7 e 0 e ;  
         r a m _ c e l l [           6 0 6 ]   =   3 2 ' h 9 c 3 7 d 6 7 5 ;  
         r a m _ c e l l [           6 0 7 ]   =   3 2 ' h b 2 7 3 6 4 8 5 ;  
         r a m _ c e l l [           6 0 8 ]   =   3 2 ' h a f 0 f e 3 f 0 ;  
         r a m _ c e l l [           6 0 9 ]   =   3 2 ' h 0 4 4 a 2 8 2 c ;  
         r a m _ c e l l [           6 1 0 ]   =   3 2 ' h 7 7 1 0 2 b 4 2 ;  
         r a m _ c e l l [           6 1 1 ]   =   3 2 ' h 9 2 a c d 2 a 4 ;  
         r a m _ c e l l [           6 1 2 ]   =   3 2 ' h b 7 f 9 5 8 d f ;  
         r a m _ c e l l [           6 1 3 ]   =   3 2 ' h 9 a f 7 b d 4 e ;  
         r a m _ c e l l [           6 1 4 ]   =   3 2 ' h 1 c 7 e 2 7 6 2 ;  
         r a m _ c e l l [           6 1 5 ]   =   3 2 ' h 1 4 b 9 7 b 4 b ;  
         r a m _ c e l l [           6 1 6 ]   =   3 2 ' h a f 8 0 e c 2 4 ;  
         r a m _ c e l l [           6 1 7 ]   =   3 2 ' h 4 a 0 6 1 d 2 5 ;  
         r a m _ c e l l [           6 1 8 ]   =   3 2 ' h c d c d 4 e d f ;  
         r a m _ c e l l [           6 1 9 ]   =   3 2 ' h 3 b e b 3 2 b a ;  
         r a m _ c e l l [           6 2 0 ]   =   3 2 ' h a 8 3 b 5 6 5 1 ;  
         r a m _ c e l l [           6 2 1 ]   =   3 2 ' h 0 e c 9 0 5 0 9 ;  
         r a m _ c e l l [           6 2 2 ]   =   3 2 ' h d c 6 b c 4 4 b ;  
         r a m _ c e l l [           6 2 3 ]   =   3 2 ' h 0 e c 5 1 0 7 e ;  
         r a m _ c e l l [           6 2 4 ]   =   3 2 ' h 6 7 e 8 0 a 2 0 ;  
         r a m _ c e l l [           6 2 5 ]   =   3 2 ' h c c 2 b 0 8 8 d ;  
         r a m _ c e l l [           6 2 6 ]   =   3 2 ' h d 8 0 e 8 b 1 5 ;  
         r a m _ c e l l [           6 2 7 ]   =   3 2 ' h f 4 e 5 8 d 2 3 ;  
         r a m _ c e l l [           6 2 8 ]   =   3 2 ' h 5 5 4 7 8 1 c c ;  
         r a m _ c e l l [           6 2 9 ]   =   3 2 ' h f d a d 6 6 b a ;  
         r a m _ c e l l [           6 3 0 ]   =   3 2 ' h c a e 0 b d 1 5 ;  
         r a m _ c e l l [           6 3 1 ]   =   3 2 ' h 6 0 9 0 5 4 f 1 ;  
         r a m _ c e l l [           6 3 2 ]   =   3 2 ' h d 7 2 7 0 2 0 9 ;  
         r a m _ c e l l [           6 3 3 ]   =   3 2 ' h 1 7 3 4 2 c c 1 ;  
         r a m _ c e l l [           6 3 4 ]   =   3 2 ' h d 8 b 9 c d 1 a ;  
         r a m _ c e l l [           6 3 5 ]   =   3 2 ' h 8 4 c f 4 8 e e ;  
         r a m _ c e l l [           6 3 6 ]   =   3 2 ' h 4 9 9 3 f f 8 4 ;  
         r a m _ c e l l [           6 3 7 ]   =   3 2 ' h 1 d c a d 0 3 8 ;  
         r a m _ c e l l [           6 3 8 ]   =   3 2 ' h 8 8 2 9 8 4 e c ;  
         r a m _ c e l l [           6 3 9 ]   =   3 2 ' h 7 f 5 8 1 a 0 2 ;  
         r a m _ c e l l [           6 4 0 ]   =   3 2 ' h d b 5 1 a 6 b 3 ;  
         r a m _ c e l l [           6 4 1 ]   =   3 2 ' h 1 b 1 e 1 b 1 9 ;  
         r a m _ c e l l [           6 4 2 ]   =   3 2 ' h 6 6 e 6 d 8 2 0 ;  
         r a m _ c e l l [           6 4 3 ]   =   3 2 ' h b 9 8 4 6 0 c f ;  
         r a m _ c e l l [           6 4 4 ]   =   3 2 ' h 7 0 5 1 3 2 7 7 ;  
         r a m _ c e l l [           6 4 5 ]   =   3 2 ' h 7 c 5 4 e 6 5 9 ;  
         r a m _ c e l l [           6 4 6 ]   =   3 2 ' h 5 8 a 4 b 3 3 8 ;  
         r a m _ c e l l [           6 4 7 ]   =   3 2 ' h e 8 8 4 d d 4 e ;  
         r a m _ c e l l [           6 4 8 ]   =   3 2 ' h 3 7 0 b a 8 9 f ;  
         r a m _ c e l l [           6 4 9 ]   =   3 2 ' h 6 a 2 2 9 f b a ;  
         r a m _ c e l l [           6 5 0 ]   =   3 2 ' h b d 9 1 4 9 a 5 ;  
         r a m _ c e l l [           6 5 1 ]   =   3 2 ' h 0 3 4 2 0 7 5 9 ;  
         r a m _ c e l l [           6 5 2 ]   =   3 2 ' h 3 c 8 b e 2 8 8 ;  
         r a m _ c e l l [           6 5 3 ]   =   3 2 ' h b 9 1 f 6 f 0 2 ;  
         r a m _ c e l l [           6 5 4 ]   =   3 2 ' h 8 a 7 7 8 8 2 c ;  
         r a m _ c e l l [           6 5 5 ]   =   3 2 ' h f f f b c 2 9 a ;  
         r a m _ c e l l [           6 5 6 ]   =   3 2 ' h 3 b c c 8 1 0 6 ;  
         r a m _ c e l l [           6 5 7 ]   =   3 2 ' h 7 5 f e 2 4 3 d ;  
         r a m _ c e l l [           6 5 8 ]   =   3 2 ' h f 3 5 7 6 9 1 3 ;  
         r a m _ c e l l [           6 5 9 ]   =   3 2 ' h c 8 f 9 5 7 5 f ;  
         r a m _ c e l l [           6 6 0 ]   =   3 2 ' h a 0 1 9 5 e e 1 ;  
         r a m _ c e l l [           6 6 1 ]   =   3 2 ' h 1 0 d 9 6 6 1 0 ;  
         r a m _ c e l l [           6 6 2 ]   =   3 2 ' h 2 2 4 6 b 2 f c ;  
         r a m _ c e l l [           6 6 3 ]   =   3 2 ' h 9 b 0 9 f 0 0 c ;  
         r a m _ c e l l [           6 6 4 ]   =   3 2 ' h a 1 1 2 7 a 5 0 ;  
         r a m _ c e l l [           6 6 5 ]   =   3 2 ' h b 7 2 f 3 e f f ;  
         r a m _ c e l l [           6 6 6 ]   =   3 2 ' h 0 b 4 8 3 4 3 c ;  
         r a m _ c e l l [           6 6 7 ]   =   3 2 ' h d 5 e 0 c 2 8 8 ;  
         r a m _ c e l l [           6 6 8 ]   =   3 2 ' h 0 4 4 e 5 9 1 a ;  
         r a m _ c e l l [           6 6 9 ]   =   3 2 ' h 2 4 5 0 3 a 9 a ;  
         r a m _ c e l l [           6 7 0 ]   =   3 2 ' h f a e c e 9 e d ;  
         r a m _ c e l l [           6 7 1 ]   =   3 2 ' h 5 3 1 9 a 9 d 2 ;  
         r a m _ c e l l [           6 7 2 ]   =   3 2 ' h e 1 f f 3 f 9 8 ;  
         r a m _ c e l l [           6 7 3 ]   =   3 2 ' h 7 8 1 d 2 e b 7 ;  
         r a m _ c e l l [           6 7 4 ]   =   3 2 ' h 9 4 7 e 1 b e 3 ;  
         r a m _ c e l l [           6 7 5 ]   =   3 2 ' h 5 c 2 9 3 0 e c ;  
         r a m _ c e l l [           6 7 6 ]   =   3 2 ' h 1 3 7 e 1 c 4 6 ;  
         r a m _ c e l l [           6 7 7 ]   =   3 2 ' h e 5 d 4 5 7 1 a ;  
         r a m _ c e l l [           6 7 8 ]   =   3 2 ' h 6 5 5 2 e 5 9 2 ;  
         r a m _ c e l l [           6 7 9 ]   =   3 2 ' h d 8 8 8 0 7 6 2 ;  
         r a m _ c e l l [           6 8 0 ]   =   3 2 ' h 6 e f a 2 e 4 5 ;  
         r a m _ c e l l [           6 8 1 ]   =   3 2 ' h 0 1 6 5 7 4 0 8 ;  
         r a m _ c e l l [           6 8 2 ]   =   3 2 ' h 5 a 0 0 9 1 6 6 ;  
         r a m _ c e l l [           6 8 3 ]   =   3 2 ' h 2 7 6 d 4 f a 2 ;  
         r a m _ c e l l [           6 8 4 ]   =   3 2 ' h 0 b 3 5 5 f a e ;  
         r a m _ c e l l [           6 8 5 ]   =   3 2 ' h e 9 6 e 3 1 e 6 ;  
         r a m _ c e l l [           6 8 6 ]   =   3 2 ' h 8 7 5 2 9 4 2 5 ;  
         r a m _ c e l l [           6 8 7 ]   =   3 2 ' h 5 9 c 6 c 9 4 b ;  
         r a m _ c e l l [           6 8 8 ]   =   3 2 ' h 1 a f 4 6 c 3 6 ;  
         r a m _ c e l l [           6 8 9 ]   =   3 2 ' h 9 7 0 0 b 5 8 f ;  
         r a m _ c e l l [           6 9 0 ]   =   3 2 ' h 8 b 5 3 d 6 b 9 ;  
         r a m _ c e l l [           6 9 1 ]   =   3 2 ' h 4 d 8 5 2 7 c a ;  
         r a m _ c e l l [           6 9 2 ]   =   3 2 ' h 6 9 3 2 c e 6 2 ;  
         r a m _ c e l l [           6 9 3 ]   =   3 2 ' h 3 c 4 9 3 d 4 1 ;  
         r a m _ c e l l [           6 9 4 ]   =   3 2 ' h b c c 7 1 b 0 f ;  
         r a m _ c e l l [           6 9 5 ]   =   3 2 ' h 9 2 5 7 8 3 e 0 ;  
         r a m _ c e l l [           6 9 6 ]   =   3 2 ' h d 7 0 2 9 3 f 7 ;  
         r a m _ c e l l [           6 9 7 ]   =   3 2 ' h d 3 2 1 f 4 c e ;  
         r a m _ c e l l [           6 9 8 ]   =   3 2 ' h c e 3 1 1 9 6 5 ;  
         r a m _ c e l l [           6 9 9 ]   =   3 2 ' h 1 c 4 4 0 4 5 2 ;  
         r a m _ c e l l [           7 0 0 ]   =   3 2 ' h 3 b 8 7 8 9 1 d ;  
         r a m _ c e l l [           7 0 1 ]   =   3 2 ' h 2 f d 5 e 8 d 5 ;  
         r a m _ c e l l [           7 0 2 ]   =   3 2 ' h 7 f 3 9 a 1 2 a ;  
         r a m _ c e l l [           7 0 3 ]   =   3 2 ' h 7 b b 8 d 5 f d ;  
         r a m _ c e l l [           7 0 4 ]   =   3 2 ' h 6 a 9 2 4 6 b 8 ;  
         r a m _ c e l l [           7 0 5 ]   =   3 2 ' h 6 5 7 7 1 8 c d ;  
         r a m _ c e l l [           7 0 6 ]   =   3 2 ' h 7 a b 1 f 6 6 3 ;  
         r a m _ c e l l [           7 0 7 ]   =   3 2 ' h e 4 b d 0 4 d 2 ;  
         r a m _ c e l l [           7 0 8 ]   =   3 2 ' h d 3 e c e 9 5 b ;  
         r a m _ c e l l [           7 0 9 ]   =   3 2 ' h e 9 4 3 2 5 1 7 ;  
         r a m _ c e l l [           7 1 0 ]   =   3 2 ' h 1 d 8 b c 9 2 2 ;  
         r a m _ c e l l [           7 1 1 ]   =   3 2 ' h e b 4 6 9 c e f ;  
         r a m _ c e l l [           7 1 2 ]   =   3 2 ' h 9 6 2 0 7 7 f c ;  
         r a m _ c e l l [           7 1 3 ]   =   3 2 ' h a 7 8 4 5 9 5 f ;  
         r a m _ c e l l [           7 1 4 ]   =   3 2 ' h d 8 f 4 7 3 3 5 ;  
         r a m _ c e l l [           7 1 5 ]   =   3 2 ' h 6 0 c 7 1 b 1 a ;  
         r a m _ c e l l [           7 1 6 ]   =   3 2 ' h 2 1 e a 5 7 7 e ;  
         r a m _ c e l l [           7 1 7 ]   =   3 2 ' h 9 a 5 d e 6 c 3 ;  
         r a m _ c e l l [           7 1 8 ]   =   3 2 ' h 5 e 1 8 5 d c 0 ;  
         r a m _ c e l l [           7 1 9 ]   =   3 2 ' h f 9 4 3 4 3 9 f ;  
         r a m _ c e l l [           7 2 0 ]   =   3 2 ' h 3 f 8 c 5 1 2 3 ;  
         r a m _ c e l l [           7 2 1 ]   =   3 2 ' h 6 c 3 6 0 6 f 7 ;  
         r a m _ c e l l [           7 2 2 ]   =   3 2 ' h 1 b 1 a 2 c 9 3 ;  
         r a m _ c e l l [           7 2 3 ]   =   3 2 ' h 6 f 6 c 3 0 f f ;  
         r a m _ c e l l [           7 2 4 ]   =   3 2 ' h 8 0 e 1 0 8 5 e ;  
         r a m _ c e l l [           7 2 5 ]   =   3 2 ' h 6 9 3 a f c a 3 ;  
         r a m _ c e l l [           7 2 6 ]   =   3 2 ' h 1 2 1 8 d b 3 1 ;  
         r a m _ c e l l [           7 2 7 ]   =   3 2 ' h a 7 2 a 2 1 f 9 ;  
         r a m _ c e l l [           7 2 8 ]   =   3 2 ' h 2 8 2 9 2 1 b 5 ;  
         r a m _ c e l l [           7 2 9 ]   =   3 2 ' h 0 b 7 0 0 0 d 0 ;  
         r a m _ c e l l [           7 3 0 ]   =   3 2 ' h 6 3 a 4 9 d 7 d ;  
         r a m _ c e l l [           7 3 1 ]   =   3 2 ' h 4 5 d 5 e 0 b 7 ;  
         r a m _ c e l l [           7 3 2 ]   =   3 2 ' h 2 c 3 f 5 4 f 9 ;  
         r a m _ c e l l [           7 3 3 ]   =   3 2 ' h a 0 9 8 9 0 0 1 ;  
         r a m _ c e l l [           7 3 4 ]   =   3 2 ' h 7 1 6 3 7 e c f ;  
         r a m _ c e l l [           7 3 5 ]   =   3 2 ' h 1 5 5 0 d 3 e 6 ;  
         r a m _ c e l l [           7 3 6 ]   =   3 2 ' h 3 f e 2 2 e d 2 ;  
         r a m _ c e l l [           7 3 7 ]   =   3 2 ' h 4 0 6 8 8 3 e 0 ;  
         r a m _ c e l l [           7 3 8 ]   =   3 2 ' h 5 5 c c 5 8 3 6 ;  
         r a m _ c e l l [           7 3 9 ]   =   3 2 ' h 7 c d d 0 8 e a ;  
         r a m _ c e l l [           7 4 0 ]   =   3 2 ' h 0 2 d 5 c 1 5 4 ;  
         r a m _ c e l l [           7 4 1 ]   =   3 2 ' h 9 d 4 7 2 a 0 a ;  
         r a m _ c e l l [           7 4 2 ]   =   3 2 ' h 2 7 b c 5 2 d 9 ;  
         r a m _ c e l l [           7 4 3 ]   =   3 2 ' h 7 e c 4 2 e 7 1 ;  
         r a m _ c e l l [           7 4 4 ]   =   3 2 ' h f d 7 3 8 5 6 a ;  
         r a m _ c e l l [           7 4 5 ]   =   3 2 ' h f 9 3 b 1 f b a ;  
         r a m _ c e l l [           7 4 6 ]   =   3 2 ' h d 8 e 9 c b 7 a ;  
         r a m _ c e l l [           7 4 7 ]   =   3 2 ' h 3 0 4 5 a d c 7 ;  
         r a m _ c e l l [           7 4 8 ]   =   3 2 ' h 4 3 5 8 c e f f ;  
         r a m _ c e l l [           7 4 9 ]   =   3 2 ' h a 6 a e 7 1 6 0 ;  
         r a m _ c e l l [           7 5 0 ]   =   3 2 ' h 0 d 3 9 5 d d a ;  
         r a m _ c e l l [           7 5 1 ]   =   3 2 ' h 5 8 a f 4 8 0 a ;  
         r a m _ c e l l [           7 5 2 ]   =   3 2 ' h 9 1 c 9 1 e 2 a ;  
         r a m _ c e l l [           7 5 3 ]   =   3 2 ' h b 9 c c e 6 1 d ;  
         r a m _ c e l l [           7 5 4 ]   =   3 2 ' h 3 1 2 d 0 5 b 1 ;  
         r a m _ c e l l [           7 5 5 ]   =   3 2 ' h 7 d 8 3 c 6 9 f ;  
         r a m _ c e l l [           7 5 6 ]   =   3 2 ' h 3 3 a b b 7 4 3 ;  
         r a m _ c e l l [           7 5 7 ]   =   3 2 ' h a e e d 0 6 8 2 ;  
         r a m _ c e l l [           7 5 8 ]   =   3 2 ' h 9 1 b f 6 c 4 f ;  
         r a m _ c e l l [           7 5 9 ]   =   3 2 ' h d 6 3 4 8 b a b ;  
         r a m _ c e l l [           7 6 0 ]   =   3 2 ' h b e d 1 3 d 2 4 ;  
         r a m _ c e l l [           7 6 1 ]   =   3 2 ' h 9 8 0 8 8 d f b ;  
         r a m _ c e l l [           7 6 2 ]   =   3 2 ' h 3 0 4 7 d d f f ;  
         r a m _ c e l l [           7 6 3 ]   =   3 2 ' h 6 7 d d 9 7 f f ;  
         r a m _ c e l l [           7 6 4 ]   =   3 2 ' h 0 e 8 c 2 d 4 4 ;  
         r a m _ c e l l [           7 6 5 ]   =   3 2 ' h 9 b 8 f f a 2 6 ;  
         r a m _ c e l l [           7 6 6 ]   =   3 2 ' h 6 e b 4 1 9 c 6 ;  
         r a m _ c e l l [           7 6 7 ]   =   3 2 ' h 5 7 6 a 1 f 6 e ;  
 e n d  
  
 e n d m o d u l e  
  
 