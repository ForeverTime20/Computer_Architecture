
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'hef2d910f;
    ram_cell[       1] = 32'h0;  // 32'hcac2afc6;
    ram_cell[       2] = 32'h0;  // 32'h37b9f3f1;
    ram_cell[       3] = 32'h0;  // 32'hdc92447c;
    ram_cell[       4] = 32'h0;  // 32'h4af5e442;
    ram_cell[       5] = 32'h0;  // 32'h9510e044;
    ram_cell[       6] = 32'h0;  // 32'hd0ea0628;
    ram_cell[       7] = 32'h0;  // 32'h0133251f;
    ram_cell[       8] = 32'h0;  // 32'hd8ba000a;
    ram_cell[       9] = 32'h0;  // 32'hb5207100;
    ram_cell[      10] = 32'h0;  // 32'h3e412433;
    ram_cell[      11] = 32'h0;  // 32'hfe9b950d;
    ram_cell[      12] = 32'h0;  // 32'h941c04cb;
    ram_cell[      13] = 32'h0;  // 32'hc0b806ad;
    ram_cell[      14] = 32'h0;  // 32'h66ec25dc;
    ram_cell[      15] = 32'h0;  // 32'h13c9457d;
    ram_cell[      16] = 32'h0;  // 32'h8d908d77;
    ram_cell[      17] = 32'h0;  // 32'hd7a4382e;
    ram_cell[      18] = 32'h0;  // 32'hf4c98001;
    ram_cell[      19] = 32'h0;  // 32'h30ab3771;
    ram_cell[      20] = 32'h0;  // 32'h19b2467a;
    ram_cell[      21] = 32'h0;  // 32'h98b1bb7c;
    ram_cell[      22] = 32'h0;  // 32'he59c2e41;
    ram_cell[      23] = 32'h0;  // 32'he01bfa89;
    ram_cell[      24] = 32'h0;  // 32'h6c58495d;
    ram_cell[      25] = 32'h0;  // 32'h7cb1f76e;
    ram_cell[      26] = 32'h0;  // 32'h368a971c;
    ram_cell[      27] = 32'h0;  // 32'ha3e5e11e;
    ram_cell[      28] = 32'h0;  // 32'h6dcf425c;
    ram_cell[      29] = 32'h0;  // 32'h254f3655;
    ram_cell[      30] = 32'h0;  // 32'h5430e0d3;
    ram_cell[      31] = 32'h0;  // 32'h232f0f15;
    ram_cell[      32] = 32'h0;  // 32'h069284f6;
    ram_cell[      33] = 32'h0;  // 32'had1add6c;
    ram_cell[      34] = 32'h0;  // 32'h05b3db72;
    ram_cell[      35] = 32'h0;  // 32'hfc0344b1;
    ram_cell[      36] = 32'h0;  // 32'hf5f62de6;
    ram_cell[      37] = 32'h0;  // 32'heaf67d3a;
    ram_cell[      38] = 32'h0;  // 32'hc6e72017;
    ram_cell[      39] = 32'h0;  // 32'h07bec8d3;
    ram_cell[      40] = 32'h0;  // 32'h32cbddcf;
    ram_cell[      41] = 32'h0;  // 32'hd8ec6106;
    ram_cell[      42] = 32'h0;  // 32'h46c2edab;
    ram_cell[      43] = 32'h0;  // 32'hf4920b93;
    ram_cell[      44] = 32'h0;  // 32'hb97548d9;
    ram_cell[      45] = 32'h0;  // 32'h691c529a;
    ram_cell[      46] = 32'h0;  // 32'h56f73615;
    ram_cell[      47] = 32'h0;  // 32'hcc033238;
    ram_cell[      48] = 32'h0;  // 32'hf6f0335d;
    ram_cell[      49] = 32'h0;  // 32'h97350f01;
    ram_cell[      50] = 32'h0;  // 32'hb45b310c;
    ram_cell[      51] = 32'h0;  // 32'h102828e9;
    ram_cell[      52] = 32'h0;  // 32'hf4a41bf6;
    ram_cell[      53] = 32'h0;  // 32'h7b220007;
    ram_cell[      54] = 32'h0;  // 32'hc9866bf0;
    ram_cell[      55] = 32'h0;  // 32'h713ead41;
    ram_cell[      56] = 32'h0;  // 32'h5a26f372;
    ram_cell[      57] = 32'h0;  // 32'hee83eed4;
    ram_cell[      58] = 32'h0;  // 32'h98221400;
    ram_cell[      59] = 32'h0;  // 32'h26635044;
    ram_cell[      60] = 32'h0;  // 32'hbeb6844e;
    ram_cell[      61] = 32'h0;  // 32'h2b7f0e7c;
    ram_cell[      62] = 32'h0;  // 32'h8243db3c;
    ram_cell[      63] = 32'h0;  // 32'h8d3c2e95;
    ram_cell[      64] = 32'h0;  // 32'h064d9d60;
    ram_cell[      65] = 32'h0;  // 32'h93a3ad2a;
    ram_cell[      66] = 32'h0;  // 32'h2502044e;
    ram_cell[      67] = 32'h0;  // 32'hec348c58;
    ram_cell[      68] = 32'h0;  // 32'h5825aaae;
    ram_cell[      69] = 32'h0;  // 32'hfb91b1fc;
    ram_cell[      70] = 32'h0;  // 32'h1859828f;
    ram_cell[      71] = 32'h0;  // 32'ha4275bda;
    ram_cell[      72] = 32'h0;  // 32'h5907b1fb;
    ram_cell[      73] = 32'h0;  // 32'h80d5e6c5;
    ram_cell[      74] = 32'h0;  // 32'h4d7646ee;
    ram_cell[      75] = 32'h0;  // 32'ha5af6d3e;
    ram_cell[      76] = 32'h0;  // 32'he4cd355c;
    ram_cell[      77] = 32'h0;  // 32'hb69d1195;
    ram_cell[      78] = 32'h0;  // 32'hdbc8e515;
    ram_cell[      79] = 32'h0;  // 32'h03387798;
    ram_cell[      80] = 32'h0;  // 32'h708b88ab;
    ram_cell[      81] = 32'h0;  // 32'h904b67af;
    ram_cell[      82] = 32'h0;  // 32'h75e87f78;
    ram_cell[      83] = 32'h0;  // 32'he40d1043;
    ram_cell[      84] = 32'h0;  // 32'h71f4f308;
    ram_cell[      85] = 32'h0;  // 32'h53b39a3d;
    ram_cell[      86] = 32'h0;  // 32'h47de073e;
    ram_cell[      87] = 32'h0;  // 32'hf6004c8e;
    ram_cell[      88] = 32'h0;  // 32'ha33e2f4d;
    ram_cell[      89] = 32'h0;  // 32'h74c4fa08;
    ram_cell[      90] = 32'h0;  // 32'ha45a5c4d;
    ram_cell[      91] = 32'h0;  // 32'he346c924;
    ram_cell[      92] = 32'h0;  // 32'h4358bd5c;
    ram_cell[      93] = 32'h0;  // 32'he7c4c037;
    ram_cell[      94] = 32'h0;  // 32'h3008f4a7;
    ram_cell[      95] = 32'h0;  // 32'h60cce51b;
    ram_cell[      96] = 32'h0;  // 32'hb2f8cd20;
    ram_cell[      97] = 32'h0;  // 32'h864236e3;
    ram_cell[      98] = 32'h0;  // 32'hfbad10d8;
    ram_cell[      99] = 32'h0;  // 32'hf49b426c;
    ram_cell[     100] = 32'h0;  // 32'h61fc5f78;
    ram_cell[     101] = 32'h0;  // 32'h48495161;
    ram_cell[     102] = 32'h0;  // 32'h0332beca;
    ram_cell[     103] = 32'h0;  // 32'hd1cc17b6;
    ram_cell[     104] = 32'h0;  // 32'h3a5c7c88;
    ram_cell[     105] = 32'h0;  // 32'h43200b9f;
    ram_cell[     106] = 32'h0;  // 32'h3711b302;
    ram_cell[     107] = 32'h0;  // 32'h0b3122b9;
    ram_cell[     108] = 32'h0;  // 32'h2a9aaac7;
    ram_cell[     109] = 32'h0;  // 32'h4a181774;
    ram_cell[     110] = 32'h0;  // 32'h2cbc185c;
    ram_cell[     111] = 32'h0;  // 32'hb86e6d2f;
    ram_cell[     112] = 32'h0;  // 32'hfe63d9e0;
    ram_cell[     113] = 32'h0;  // 32'hce840f80;
    ram_cell[     114] = 32'h0;  // 32'h3f5ced79;
    ram_cell[     115] = 32'h0;  // 32'h58588eb8;
    ram_cell[     116] = 32'h0;  // 32'hdccab3a6;
    ram_cell[     117] = 32'h0;  // 32'h2694c2b8;
    ram_cell[     118] = 32'h0;  // 32'h8429e656;
    ram_cell[     119] = 32'h0;  // 32'h30ba8adc;
    ram_cell[     120] = 32'h0;  // 32'hd2319b6e;
    ram_cell[     121] = 32'h0;  // 32'ha061eb6b;
    ram_cell[     122] = 32'h0;  // 32'h1421f7c8;
    ram_cell[     123] = 32'h0;  // 32'h0f209e4d;
    ram_cell[     124] = 32'h0;  // 32'hdb3a9389;
    ram_cell[     125] = 32'h0;  // 32'hacfffd76;
    ram_cell[     126] = 32'h0;  // 32'h49019103;
    ram_cell[     127] = 32'h0;  // 32'h304d6210;
    ram_cell[     128] = 32'h0;  // 32'hf2f003df;
    ram_cell[     129] = 32'h0;  // 32'h4384628e;
    ram_cell[     130] = 32'h0;  // 32'hbd5dc668;
    ram_cell[     131] = 32'h0;  // 32'h20a7a4cb;
    ram_cell[     132] = 32'h0;  // 32'hbe7de225;
    ram_cell[     133] = 32'h0;  // 32'h3a3c73cd;
    ram_cell[     134] = 32'h0;  // 32'h8439a659;
    ram_cell[     135] = 32'h0;  // 32'hdfe6275e;
    ram_cell[     136] = 32'h0;  // 32'h1e21d413;
    ram_cell[     137] = 32'h0;  // 32'h43d6b1df;
    ram_cell[     138] = 32'h0;  // 32'hc46a06ed;
    ram_cell[     139] = 32'h0;  // 32'ha91db16c;
    ram_cell[     140] = 32'h0;  // 32'h27733819;
    ram_cell[     141] = 32'h0;  // 32'he73a4a52;
    ram_cell[     142] = 32'h0;  // 32'hf8dcd530;
    ram_cell[     143] = 32'h0;  // 32'h63f70fa9;
    ram_cell[     144] = 32'h0;  // 32'hb23b9941;
    ram_cell[     145] = 32'h0;  // 32'hed157b62;
    ram_cell[     146] = 32'h0;  // 32'h3c9c553f;
    ram_cell[     147] = 32'h0;  // 32'hd0964663;
    ram_cell[     148] = 32'h0;  // 32'h80709f77;
    ram_cell[     149] = 32'h0;  // 32'h7a8ac36b;
    ram_cell[     150] = 32'h0;  // 32'hc41d4e9b;
    ram_cell[     151] = 32'h0;  // 32'hfdcd5dd1;
    ram_cell[     152] = 32'h0;  // 32'hdf2dc9f8;
    ram_cell[     153] = 32'h0;  // 32'hfe413582;
    ram_cell[     154] = 32'h0;  // 32'h2bc5d186;
    ram_cell[     155] = 32'h0;  // 32'h3869a465;
    ram_cell[     156] = 32'h0;  // 32'h9991cc69;
    ram_cell[     157] = 32'h0;  // 32'h0b020951;
    ram_cell[     158] = 32'h0;  // 32'h2edc7ad4;
    ram_cell[     159] = 32'h0;  // 32'haed1c13b;
    ram_cell[     160] = 32'h0;  // 32'h8c1aa012;
    ram_cell[     161] = 32'h0;  // 32'h9db426e2;
    ram_cell[     162] = 32'h0;  // 32'h85b50ab2;
    ram_cell[     163] = 32'h0;  // 32'h2586c533;
    ram_cell[     164] = 32'h0;  // 32'h19af9d00;
    ram_cell[     165] = 32'h0;  // 32'hd3795976;
    ram_cell[     166] = 32'h0;  // 32'hc56d8f7b;
    ram_cell[     167] = 32'h0;  // 32'h7a1fa280;
    ram_cell[     168] = 32'h0;  // 32'h0beaad5f;
    ram_cell[     169] = 32'h0;  // 32'h9dfdd518;
    ram_cell[     170] = 32'h0;  // 32'hf0f3f578;
    ram_cell[     171] = 32'h0;  // 32'h111dfdf8;
    ram_cell[     172] = 32'h0;  // 32'hc861e967;
    ram_cell[     173] = 32'h0;  // 32'h543a3fdd;
    ram_cell[     174] = 32'h0;  // 32'haf1d759d;
    ram_cell[     175] = 32'h0;  // 32'h5b910529;
    ram_cell[     176] = 32'h0;  // 32'h7549c395;
    ram_cell[     177] = 32'h0;  // 32'h828664b8;
    ram_cell[     178] = 32'h0;  // 32'h54ee8b76;
    ram_cell[     179] = 32'h0;  // 32'had9157d6;
    ram_cell[     180] = 32'h0;  // 32'h2c10a3a5;
    ram_cell[     181] = 32'h0;  // 32'haec8475e;
    ram_cell[     182] = 32'h0;  // 32'h33e58ca3;
    ram_cell[     183] = 32'h0;  // 32'hc48a4269;
    ram_cell[     184] = 32'h0;  // 32'ha8cea106;
    ram_cell[     185] = 32'h0;  // 32'h296e7477;
    ram_cell[     186] = 32'h0;  // 32'h7936649f;
    ram_cell[     187] = 32'h0;  // 32'h9a7082e4;
    ram_cell[     188] = 32'h0;  // 32'h8647c471;
    ram_cell[     189] = 32'h0;  // 32'hd723b705;
    ram_cell[     190] = 32'h0;  // 32'h4944454d;
    ram_cell[     191] = 32'h0;  // 32'haf1b362e;
    ram_cell[     192] = 32'h0;  // 32'hf2b11e7c;
    ram_cell[     193] = 32'h0;  // 32'h1ab72c37;
    ram_cell[     194] = 32'h0;  // 32'hf70f8477;
    ram_cell[     195] = 32'h0;  // 32'h8add12f2;
    ram_cell[     196] = 32'h0;  // 32'h2ebf7010;
    ram_cell[     197] = 32'h0;  // 32'hb06a6a1f;
    ram_cell[     198] = 32'h0;  // 32'h9f16b5ac;
    ram_cell[     199] = 32'h0;  // 32'h17638cc5;
    ram_cell[     200] = 32'h0;  // 32'h4e7165eb;
    ram_cell[     201] = 32'h0;  // 32'hc240829d;
    ram_cell[     202] = 32'h0;  // 32'h5d0c869e;
    ram_cell[     203] = 32'h0;  // 32'hefaa5566;
    ram_cell[     204] = 32'h0;  // 32'h872d7f0f;
    ram_cell[     205] = 32'h0;  // 32'h6ab7d1a9;
    ram_cell[     206] = 32'h0;  // 32'hb3c3a376;
    ram_cell[     207] = 32'h0;  // 32'he73cc1b3;
    ram_cell[     208] = 32'h0;  // 32'ha4a306b2;
    ram_cell[     209] = 32'h0;  // 32'hbeb15104;
    ram_cell[     210] = 32'h0;  // 32'he70d3981;
    ram_cell[     211] = 32'h0;  // 32'h70daca48;
    ram_cell[     212] = 32'h0;  // 32'h08dd62e3;
    ram_cell[     213] = 32'h0;  // 32'ha6697ece;
    ram_cell[     214] = 32'h0;  // 32'h068f3aa3;
    ram_cell[     215] = 32'h0;  // 32'h03219e61;
    ram_cell[     216] = 32'h0;  // 32'hdf3e7629;
    ram_cell[     217] = 32'h0;  // 32'hbd252939;
    ram_cell[     218] = 32'h0;  // 32'h7d412e33;
    ram_cell[     219] = 32'h0;  // 32'h9b832ac6;
    ram_cell[     220] = 32'h0;  // 32'h0aa05de6;
    ram_cell[     221] = 32'h0;  // 32'h7a99b0a2;
    ram_cell[     222] = 32'h0;  // 32'h108deb5c;
    ram_cell[     223] = 32'h0;  // 32'hb97e4180;
    ram_cell[     224] = 32'h0;  // 32'hac7fe810;
    ram_cell[     225] = 32'h0;  // 32'h9536e3db;
    ram_cell[     226] = 32'h0;  // 32'hc6340613;
    ram_cell[     227] = 32'h0;  // 32'h820688db;
    ram_cell[     228] = 32'h0;  // 32'hedb9303b;
    ram_cell[     229] = 32'h0;  // 32'h9fe4cb8e;
    ram_cell[     230] = 32'h0;  // 32'h3c1349f5;
    ram_cell[     231] = 32'h0;  // 32'h19f60640;
    ram_cell[     232] = 32'h0;  // 32'hb103a4a7;
    ram_cell[     233] = 32'h0;  // 32'h29b42cc8;
    ram_cell[     234] = 32'h0;  // 32'hc5835177;
    ram_cell[     235] = 32'h0;  // 32'h22937328;
    ram_cell[     236] = 32'h0;  // 32'h0337a0de;
    ram_cell[     237] = 32'h0;  // 32'h6317747f;
    ram_cell[     238] = 32'h0;  // 32'hafd8b7f0;
    ram_cell[     239] = 32'h0;  // 32'h378a8eb7;
    ram_cell[     240] = 32'h0;  // 32'hc68484a8;
    ram_cell[     241] = 32'h0;  // 32'h833ca399;
    ram_cell[     242] = 32'h0;  // 32'h452b8a34;
    ram_cell[     243] = 32'h0;  // 32'h079ed023;
    ram_cell[     244] = 32'h0;  // 32'h9e3b1da4;
    ram_cell[     245] = 32'h0;  // 32'hd4f32555;
    ram_cell[     246] = 32'h0;  // 32'hdf6b2168;
    ram_cell[     247] = 32'h0;  // 32'h8da4a3c0;
    ram_cell[     248] = 32'h0;  // 32'hf2ef828b;
    ram_cell[     249] = 32'h0;  // 32'h0c8ee6a4;
    ram_cell[     250] = 32'h0;  // 32'h31ae0849;
    ram_cell[     251] = 32'h0;  // 32'h9f0356b7;
    ram_cell[     252] = 32'h0;  // 32'h254ce6c4;
    ram_cell[     253] = 32'h0;  // 32'h60b817e7;
    ram_cell[     254] = 32'h0;  // 32'h1c33b98c;
    ram_cell[     255] = 32'h0;  // 32'h2d64e6e5;
    // src matrix A
    ram_cell[     256] = 32'hc3bbcca6;
    ram_cell[     257] = 32'hd6224481;
    ram_cell[     258] = 32'he57924af;
    ram_cell[     259] = 32'h2dd8fcfc;
    ram_cell[     260] = 32'h9e4f7c11;
    ram_cell[     261] = 32'h8755911e;
    ram_cell[     262] = 32'hcb5665aa;
    ram_cell[     263] = 32'ha6bd8f33;
    ram_cell[     264] = 32'h35410441;
    ram_cell[     265] = 32'h425d2d68;
    ram_cell[     266] = 32'hf44ac70e;
    ram_cell[     267] = 32'h0d86e121;
    ram_cell[     268] = 32'h5e97196a;
    ram_cell[     269] = 32'hcd4bf0e5;
    ram_cell[     270] = 32'h0d627792;
    ram_cell[     271] = 32'hb75f2d3d;
    ram_cell[     272] = 32'h84e265d0;
    ram_cell[     273] = 32'h722e6b37;
    ram_cell[     274] = 32'ha3a8e8f1;
    ram_cell[     275] = 32'h5e5f2a09;
    ram_cell[     276] = 32'h9d783304;
    ram_cell[     277] = 32'hb082b07e;
    ram_cell[     278] = 32'h08cd00ca;
    ram_cell[     279] = 32'hda0f515d;
    ram_cell[     280] = 32'hbc64ea71;
    ram_cell[     281] = 32'h43d4fca9;
    ram_cell[     282] = 32'h9196fc16;
    ram_cell[     283] = 32'hd4cf46e5;
    ram_cell[     284] = 32'h32cd89d5;
    ram_cell[     285] = 32'h936de192;
    ram_cell[     286] = 32'h152d3640;
    ram_cell[     287] = 32'h5c54d2b1;
    ram_cell[     288] = 32'h41a72345;
    ram_cell[     289] = 32'h055b25d2;
    ram_cell[     290] = 32'h959d570a;
    ram_cell[     291] = 32'h5f190d74;
    ram_cell[     292] = 32'h78fa8603;
    ram_cell[     293] = 32'h5e691a6b;
    ram_cell[     294] = 32'h9fc6b162;
    ram_cell[     295] = 32'he430fd23;
    ram_cell[     296] = 32'h9ea768c8;
    ram_cell[     297] = 32'h2f5d233e;
    ram_cell[     298] = 32'h619deea3;
    ram_cell[     299] = 32'h335698a2;
    ram_cell[     300] = 32'hacde6fc7;
    ram_cell[     301] = 32'h80880700;
    ram_cell[     302] = 32'hf2c23485;
    ram_cell[     303] = 32'h69a3e84d;
    ram_cell[     304] = 32'h55e89669;
    ram_cell[     305] = 32'h919155f2;
    ram_cell[     306] = 32'hc9b09ad9;
    ram_cell[     307] = 32'h612f3c90;
    ram_cell[     308] = 32'hd4e526f8;
    ram_cell[     309] = 32'h3189c638;
    ram_cell[     310] = 32'he35b0656;
    ram_cell[     311] = 32'hd6e14882;
    ram_cell[     312] = 32'hf707309a;
    ram_cell[     313] = 32'h0bd9bc1f;
    ram_cell[     314] = 32'ha4522b9f;
    ram_cell[     315] = 32'h5d614934;
    ram_cell[     316] = 32'hd27562c7;
    ram_cell[     317] = 32'h51ac7084;
    ram_cell[     318] = 32'hbd7c106a;
    ram_cell[     319] = 32'hfcf40b5d;
    ram_cell[     320] = 32'h4459fe44;
    ram_cell[     321] = 32'h44ed3762;
    ram_cell[     322] = 32'hc5523a88;
    ram_cell[     323] = 32'h4284976c;
    ram_cell[     324] = 32'ha1f4c7da;
    ram_cell[     325] = 32'hd261302f;
    ram_cell[     326] = 32'h64faaa0d;
    ram_cell[     327] = 32'hbfcbd2ce;
    ram_cell[     328] = 32'he6c095e2;
    ram_cell[     329] = 32'h865bbc8f;
    ram_cell[     330] = 32'hefeccbec;
    ram_cell[     331] = 32'hae6617c6;
    ram_cell[     332] = 32'h8ba1dedc;
    ram_cell[     333] = 32'he51966df;
    ram_cell[     334] = 32'h1a48e0f2;
    ram_cell[     335] = 32'h0b85a996;
    ram_cell[     336] = 32'h2ce6d40f;
    ram_cell[     337] = 32'ha4266e38;
    ram_cell[     338] = 32'h6a17f2c9;
    ram_cell[     339] = 32'hba5daadd;
    ram_cell[     340] = 32'h6b55bc03;
    ram_cell[     341] = 32'h68c9f6d5;
    ram_cell[     342] = 32'h869e3459;
    ram_cell[     343] = 32'h7a78b7eb;
    ram_cell[     344] = 32'hcecfebae;
    ram_cell[     345] = 32'haadf002f;
    ram_cell[     346] = 32'h2c831d1e;
    ram_cell[     347] = 32'h51793619;
    ram_cell[     348] = 32'hcf979faf;
    ram_cell[     349] = 32'h71363370;
    ram_cell[     350] = 32'hc0bcd98a;
    ram_cell[     351] = 32'h86cc0c4e;
    ram_cell[     352] = 32'h84f9c22c;
    ram_cell[     353] = 32'h2b3f08cb;
    ram_cell[     354] = 32'hd8d6ad4f;
    ram_cell[     355] = 32'h5057f3bf;
    ram_cell[     356] = 32'hf3dec8d0;
    ram_cell[     357] = 32'h861bfc1a;
    ram_cell[     358] = 32'ha86c1e8c;
    ram_cell[     359] = 32'h29c6f622;
    ram_cell[     360] = 32'hd4fa13a4;
    ram_cell[     361] = 32'ha768ec84;
    ram_cell[     362] = 32'h65f9d036;
    ram_cell[     363] = 32'hd81d65c6;
    ram_cell[     364] = 32'hfc494811;
    ram_cell[     365] = 32'h5d27eff2;
    ram_cell[     366] = 32'h92103b79;
    ram_cell[     367] = 32'h9b5bf7c3;
    ram_cell[     368] = 32'ha5ff9a89;
    ram_cell[     369] = 32'h84e6c357;
    ram_cell[     370] = 32'h0d0f536e;
    ram_cell[     371] = 32'h04a046ea;
    ram_cell[     372] = 32'h2051a78e;
    ram_cell[     373] = 32'h426a0e94;
    ram_cell[     374] = 32'h292ad71e;
    ram_cell[     375] = 32'ha0ff6a0e;
    ram_cell[     376] = 32'h6d1432d1;
    ram_cell[     377] = 32'hbbbdbb22;
    ram_cell[     378] = 32'h56010493;
    ram_cell[     379] = 32'hed9d0be6;
    ram_cell[     380] = 32'h67664cd8;
    ram_cell[     381] = 32'h39306bc1;
    ram_cell[     382] = 32'h8aefdccc;
    ram_cell[     383] = 32'h8130fb5c;
    ram_cell[     384] = 32'hac956fa6;
    ram_cell[     385] = 32'h052e4628;
    ram_cell[     386] = 32'haa4a2e41;
    ram_cell[     387] = 32'h3f7b2c81;
    ram_cell[     388] = 32'h83e8dc7d;
    ram_cell[     389] = 32'h03b90878;
    ram_cell[     390] = 32'h6d55bf15;
    ram_cell[     391] = 32'hd26bc15b;
    ram_cell[     392] = 32'hbbe96ee8;
    ram_cell[     393] = 32'ha4fa28f3;
    ram_cell[     394] = 32'ha494a97c;
    ram_cell[     395] = 32'h87a04455;
    ram_cell[     396] = 32'h6cd65d10;
    ram_cell[     397] = 32'h9946aab5;
    ram_cell[     398] = 32'h0d97ab00;
    ram_cell[     399] = 32'h2f92360d;
    ram_cell[     400] = 32'h956ebdf3;
    ram_cell[     401] = 32'h4d6dd3fc;
    ram_cell[     402] = 32'h5a42add0;
    ram_cell[     403] = 32'hfa222b53;
    ram_cell[     404] = 32'ha89f5013;
    ram_cell[     405] = 32'he899f84d;
    ram_cell[     406] = 32'h2c68b76a;
    ram_cell[     407] = 32'hb2563c0e;
    ram_cell[     408] = 32'h9b5c4ef3;
    ram_cell[     409] = 32'hd336c45d;
    ram_cell[     410] = 32'h22b6a593;
    ram_cell[     411] = 32'h628e713b;
    ram_cell[     412] = 32'heffd7aa5;
    ram_cell[     413] = 32'he0dc4dfb;
    ram_cell[     414] = 32'hc37725ed;
    ram_cell[     415] = 32'h5e0253f1;
    ram_cell[     416] = 32'h7df6671e;
    ram_cell[     417] = 32'he1ae024c;
    ram_cell[     418] = 32'he1245ff1;
    ram_cell[     419] = 32'h48620017;
    ram_cell[     420] = 32'h067f62e4;
    ram_cell[     421] = 32'hef8c6bf5;
    ram_cell[     422] = 32'hc6cc5a2b;
    ram_cell[     423] = 32'hea654932;
    ram_cell[     424] = 32'h2baa8795;
    ram_cell[     425] = 32'h6829716e;
    ram_cell[     426] = 32'h7fa972e5;
    ram_cell[     427] = 32'hff707104;
    ram_cell[     428] = 32'h3a1c0446;
    ram_cell[     429] = 32'hb8747754;
    ram_cell[     430] = 32'h07a39938;
    ram_cell[     431] = 32'h1610b6fe;
    ram_cell[     432] = 32'h479531c5;
    ram_cell[     433] = 32'h957643eb;
    ram_cell[     434] = 32'he89e1bba;
    ram_cell[     435] = 32'h4ac4ae86;
    ram_cell[     436] = 32'hd21dd927;
    ram_cell[     437] = 32'h10d50e71;
    ram_cell[     438] = 32'hf8642a71;
    ram_cell[     439] = 32'hd1ad56a8;
    ram_cell[     440] = 32'h15874c98;
    ram_cell[     441] = 32'hb00a806c;
    ram_cell[     442] = 32'h2a5ec322;
    ram_cell[     443] = 32'h41f87192;
    ram_cell[     444] = 32'haec30d74;
    ram_cell[     445] = 32'h66d93e4f;
    ram_cell[     446] = 32'hd5adb554;
    ram_cell[     447] = 32'h5122ff6b;
    ram_cell[     448] = 32'h181ca871;
    ram_cell[     449] = 32'h272af914;
    ram_cell[     450] = 32'h6fefd9fd;
    ram_cell[     451] = 32'hfa225b3f;
    ram_cell[     452] = 32'h97151e47;
    ram_cell[     453] = 32'hd4cd6ddb;
    ram_cell[     454] = 32'h31b80a0a;
    ram_cell[     455] = 32'haabba76e;
    ram_cell[     456] = 32'h005ee68a;
    ram_cell[     457] = 32'hb1339cad;
    ram_cell[     458] = 32'hf6844be8;
    ram_cell[     459] = 32'h447ed3b7;
    ram_cell[     460] = 32'h1c9a4545;
    ram_cell[     461] = 32'hab1693d9;
    ram_cell[     462] = 32'h3eee12e0;
    ram_cell[     463] = 32'h51d481d9;
    ram_cell[     464] = 32'h084fb282;
    ram_cell[     465] = 32'hc60b0647;
    ram_cell[     466] = 32'h6d569ad1;
    ram_cell[     467] = 32'hd29fecd9;
    ram_cell[     468] = 32'h842ef4c9;
    ram_cell[     469] = 32'hd6c8c4e9;
    ram_cell[     470] = 32'h02a241cd;
    ram_cell[     471] = 32'hcf04d242;
    ram_cell[     472] = 32'h797446b6;
    ram_cell[     473] = 32'hc73a0687;
    ram_cell[     474] = 32'h1c56b739;
    ram_cell[     475] = 32'he85230f9;
    ram_cell[     476] = 32'h516f71fd;
    ram_cell[     477] = 32'haf3b82d4;
    ram_cell[     478] = 32'hc7275c32;
    ram_cell[     479] = 32'h2a528225;
    ram_cell[     480] = 32'hcd0e193f;
    ram_cell[     481] = 32'hd9cf312f;
    ram_cell[     482] = 32'hb4ac04d5;
    ram_cell[     483] = 32'h5f8f6dfe;
    ram_cell[     484] = 32'hda0f0f7e;
    ram_cell[     485] = 32'h8f0ae556;
    ram_cell[     486] = 32'h88632fc4;
    ram_cell[     487] = 32'hbe09b61c;
    ram_cell[     488] = 32'hb9abfc2d;
    ram_cell[     489] = 32'h98af2a42;
    ram_cell[     490] = 32'h3f096cc2;
    ram_cell[     491] = 32'h40ef5af1;
    ram_cell[     492] = 32'hb40761f7;
    ram_cell[     493] = 32'hc873481d;
    ram_cell[     494] = 32'h7a4d337f;
    ram_cell[     495] = 32'h6e509138;
    ram_cell[     496] = 32'hf6045571;
    ram_cell[     497] = 32'heaf9c1a7;
    ram_cell[     498] = 32'h4a8c58f9;
    ram_cell[     499] = 32'hc44e54ca;
    ram_cell[     500] = 32'h76b379d3;
    ram_cell[     501] = 32'h96a1fd94;
    ram_cell[     502] = 32'he5c30308;
    ram_cell[     503] = 32'h35bba4b9;
    ram_cell[     504] = 32'h33ba7cde;
    ram_cell[     505] = 32'h5e865d26;
    ram_cell[     506] = 32'he6f844c8;
    ram_cell[     507] = 32'hf5c8fa91;
    ram_cell[     508] = 32'h9d6069ac;
    ram_cell[     509] = 32'h17fa127e;
    ram_cell[     510] = 32'hc53e7561;
    ram_cell[     511] = 32'hd78037f3;
    // src matrix B
    ram_cell[     512] = 32'h08c3831e;
    ram_cell[     513] = 32'h93694116;
    ram_cell[     514] = 32'h8835ce6f;
    ram_cell[     515] = 32'h265dcab7;
    ram_cell[     516] = 32'hdae194d0;
    ram_cell[     517] = 32'h59b9ef0c;
    ram_cell[     518] = 32'hd4af98c6;
    ram_cell[     519] = 32'hf47a143e;
    ram_cell[     520] = 32'h91544bff;
    ram_cell[     521] = 32'he482bb8f;
    ram_cell[     522] = 32'h7a3a22e3;
    ram_cell[     523] = 32'h5d2f902e;
    ram_cell[     524] = 32'ha7a7cbe1;
    ram_cell[     525] = 32'hebbbe686;
    ram_cell[     526] = 32'h21a10558;
    ram_cell[     527] = 32'hf99c37c6;
    ram_cell[     528] = 32'hdaaf7d70;
    ram_cell[     529] = 32'hb72198ee;
    ram_cell[     530] = 32'h60afbce5;
    ram_cell[     531] = 32'hedbbf8fa;
    ram_cell[     532] = 32'hd2cffbee;
    ram_cell[     533] = 32'h1335d033;
    ram_cell[     534] = 32'h3b89d1ee;
    ram_cell[     535] = 32'hbb3f7f61;
    ram_cell[     536] = 32'h63acb695;
    ram_cell[     537] = 32'hfabee023;
    ram_cell[     538] = 32'ha10a187a;
    ram_cell[     539] = 32'h8764571a;
    ram_cell[     540] = 32'h7c39b916;
    ram_cell[     541] = 32'h743b19d4;
    ram_cell[     542] = 32'hfbda278c;
    ram_cell[     543] = 32'h1bbca223;
    ram_cell[     544] = 32'hf96ebbc0;
    ram_cell[     545] = 32'h7a552683;
    ram_cell[     546] = 32'h92f86df0;
    ram_cell[     547] = 32'h7a7a0993;
    ram_cell[     548] = 32'had1369fe;
    ram_cell[     549] = 32'hc0114668;
    ram_cell[     550] = 32'h886497ee;
    ram_cell[     551] = 32'hd586f633;
    ram_cell[     552] = 32'h31d84d5a;
    ram_cell[     553] = 32'h3ce8b037;
    ram_cell[     554] = 32'h13d87188;
    ram_cell[     555] = 32'h3c8f7177;
    ram_cell[     556] = 32'h684f3bcd;
    ram_cell[     557] = 32'h34c3b692;
    ram_cell[     558] = 32'hd55415e0;
    ram_cell[     559] = 32'hd665dc9a;
    ram_cell[     560] = 32'h28748887;
    ram_cell[     561] = 32'h522c83d3;
    ram_cell[     562] = 32'h8d5258af;
    ram_cell[     563] = 32'h31bc4bf0;
    ram_cell[     564] = 32'hc499da68;
    ram_cell[     565] = 32'h0aae697d;
    ram_cell[     566] = 32'he6a6a782;
    ram_cell[     567] = 32'h3ded9a49;
    ram_cell[     568] = 32'hcb16e9b7;
    ram_cell[     569] = 32'h9909c5a2;
    ram_cell[     570] = 32'hf6647d76;
    ram_cell[     571] = 32'h8feb9bf0;
    ram_cell[     572] = 32'h395167a2;
    ram_cell[     573] = 32'h753b92b0;
    ram_cell[     574] = 32'h25507db1;
    ram_cell[     575] = 32'h695004f8;
    ram_cell[     576] = 32'ha6aa6d96;
    ram_cell[     577] = 32'h68be610c;
    ram_cell[     578] = 32'ha6e51476;
    ram_cell[     579] = 32'h1ddd8afb;
    ram_cell[     580] = 32'hcae42ab8;
    ram_cell[     581] = 32'h2b50a6d3;
    ram_cell[     582] = 32'ha034f3a9;
    ram_cell[     583] = 32'h1279453e;
    ram_cell[     584] = 32'h39e169f1;
    ram_cell[     585] = 32'h5f2f498e;
    ram_cell[     586] = 32'hff34dea4;
    ram_cell[     587] = 32'h78cfd9f7;
    ram_cell[     588] = 32'heb7fa21b;
    ram_cell[     589] = 32'h11b6b027;
    ram_cell[     590] = 32'hd6886276;
    ram_cell[     591] = 32'h029fc205;
    ram_cell[     592] = 32'h97fe74a8;
    ram_cell[     593] = 32'ha1b71224;
    ram_cell[     594] = 32'h5390703c;
    ram_cell[     595] = 32'hc391129d;
    ram_cell[     596] = 32'hc4440ffa;
    ram_cell[     597] = 32'h35edb57c;
    ram_cell[     598] = 32'he471744e;
    ram_cell[     599] = 32'h75121591;
    ram_cell[     600] = 32'hfd5a2462;
    ram_cell[     601] = 32'hb01ae8c6;
    ram_cell[     602] = 32'h89498586;
    ram_cell[     603] = 32'h9c9f90fb;
    ram_cell[     604] = 32'he185524f;
    ram_cell[     605] = 32'he03fbef7;
    ram_cell[     606] = 32'h48e288b3;
    ram_cell[     607] = 32'h9850f855;
    ram_cell[     608] = 32'h80462cf6;
    ram_cell[     609] = 32'h51dbefb4;
    ram_cell[     610] = 32'hfe438fe4;
    ram_cell[     611] = 32'h91349c0d;
    ram_cell[     612] = 32'h7b540ecc;
    ram_cell[     613] = 32'h20bd9463;
    ram_cell[     614] = 32'h8640c0d0;
    ram_cell[     615] = 32'h9d27b917;
    ram_cell[     616] = 32'h779f74a1;
    ram_cell[     617] = 32'ha82fe701;
    ram_cell[     618] = 32'hf2068a17;
    ram_cell[     619] = 32'h72c83f6c;
    ram_cell[     620] = 32'hf1dbbd9b;
    ram_cell[     621] = 32'h810ef8ab;
    ram_cell[     622] = 32'ha8aeab30;
    ram_cell[     623] = 32'hf2014f1c;
    ram_cell[     624] = 32'h696f8310;
    ram_cell[     625] = 32'h7ac14e34;
    ram_cell[     626] = 32'ha105ecdf;
    ram_cell[     627] = 32'h6307474c;
    ram_cell[     628] = 32'hf3809b9d;
    ram_cell[     629] = 32'h0890c67a;
    ram_cell[     630] = 32'hd0b582b2;
    ram_cell[     631] = 32'hb58daa56;
    ram_cell[     632] = 32'h36dfd6c7;
    ram_cell[     633] = 32'h2f492b16;
    ram_cell[     634] = 32'h3be2f073;
    ram_cell[     635] = 32'hb0ebad52;
    ram_cell[     636] = 32'hccc839ad;
    ram_cell[     637] = 32'hcc7fb6c7;
    ram_cell[     638] = 32'h13070213;
    ram_cell[     639] = 32'h36114b89;
    ram_cell[     640] = 32'h6be9d3c4;
    ram_cell[     641] = 32'h4a1802d7;
    ram_cell[     642] = 32'h71429d39;
    ram_cell[     643] = 32'hbcef2013;
    ram_cell[     644] = 32'h446566ab;
    ram_cell[     645] = 32'h9440ab92;
    ram_cell[     646] = 32'h2bc96475;
    ram_cell[     647] = 32'ha72987bf;
    ram_cell[     648] = 32'h23e55789;
    ram_cell[     649] = 32'h28f7ab2e;
    ram_cell[     650] = 32'hb769a1ce;
    ram_cell[     651] = 32'hf0393bd1;
    ram_cell[     652] = 32'h8fdc9789;
    ram_cell[     653] = 32'h92d6594c;
    ram_cell[     654] = 32'hcffc82dd;
    ram_cell[     655] = 32'h5f853fe3;
    ram_cell[     656] = 32'hd5e487bb;
    ram_cell[     657] = 32'h13eb8a26;
    ram_cell[     658] = 32'hb9671482;
    ram_cell[     659] = 32'h8ef137c7;
    ram_cell[     660] = 32'h775596de;
    ram_cell[     661] = 32'h5b60a25e;
    ram_cell[     662] = 32'h94f5af96;
    ram_cell[     663] = 32'h162e036d;
    ram_cell[     664] = 32'h4ffbdb25;
    ram_cell[     665] = 32'h33bba62b;
    ram_cell[     666] = 32'h5cb78aa9;
    ram_cell[     667] = 32'h3f44cfcc;
    ram_cell[     668] = 32'h837db818;
    ram_cell[     669] = 32'h373d9f34;
    ram_cell[     670] = 32'h37714bdc;
    ram_cell[     671] = 32'h7bf421ac;
    ram_cell[     672] = 32'h5bb1a9f5;
    ram_cell[     673] = 32'h489a30a7;
    ram_cell[     674] = 32'h210e34e0;
    ram_cell[     675] = 32'h01d28e5f;
    ram_cell[     676] = 32'h7be00ec1;
    ram_cell[     677] = 32'h555d19ae;
    ram_cell[     678] = 32'hf392de1c;
    ram_cell[     679] = 32'hb5fd9adf;
    ram_cell[     680] = 32'hb574e656;
    ram_cell[     681] = 32'h79a8fa7a;
    ram_cell[     682] = 32'h4cea333b;
    ram_cell[     683] = 32'hda302e8d;
    ram_cell[     684] = 32'hb9148ae9;
    ram_cell[     685] = 32'h5ac487e9;
    ram_cell[     686] = 32'he1c19d64;
    ram_cell[     687] = 32'h3d392fa3;
    ram_cell[     688] = 32'hc58a1036;
    ram_cell[     689] = 32'h9d9db370;
    ram_cell[     690] = 32'ha13c1a9a;
    ram_cell[     691] = 32'h0bc29d5b;
    ram_cell[     692] = 32'h0a97d9a3;
    ram_cell[     693] = 32'h2dd5832f;
    ram_cell[     694] = 32'he0014446;
    ram_cell[     695] = 32'h7f77754a;
    ram_cell[     696] = 32'h69068906;
    ram_cell[     697] = 32'h5a796012;
    ram_cell[     698] = 32'h0fb19261;
    ram_cell[     699] = 32'hb6bbfe26;
    ram_cell[     700] = 32'hb7a827ae;
    ram_cell[     701] = 32'h4be235a5;
    ram_cell[     702] = 32'hf6b9255e;
    ram_cell[     703] = 32'h6c4fb772;
    ram_cell[     704] = 32'h638eae25;
    ram_cell[     705] = 32'hc347785b;
    ram_cell[     706] = 32'h2948ebf7;
    ram_cell[     707] = 32'hd8245334;
    ram_cell[     708] = 32'hcbdc6e18;
    ram_cell[     709] = 32'h26212617;
    ram_cell[     710] = 32'h6247c381;
    ram_cell[     711] = 32'h4f489a13;
    ram_cell[     712] = 32'he7b25351;
    ram_cell[     713] = 32'h8f2378c0;
    ram_cell[     714] = 32'h75648410;
    ram_cell[     715] = 32'h488c408b;
    ram_cell[     716] = 32'hb65e7eb8;
    ram_cell[     717] = 32'hcc7d366a;
    ram_cell[     718] = 32'h0df97f7e;
    ram_cell[     719] = 32'ha88cff3c;
    ram_cell[     720] = 32'hf13b559b;
    ram_cell[     721] = 32'h4af4fd26;
    ram_cell[     722] = 32'hadc9a824;
    ram_cell[     723] = 32'hbbb25211;
    ram_cell[     724] = 32'h6ead7de2;
    ram_cell[     725] = 32'h911b2a6f;
    ram_cell[     726] = 32'hfe93864f;
    ram_cell[     727] = 32'h1c7cb4a7;
    ram_cell[     728] = 32'hd92baecb;
    ram_cell[     729] = 32'he1ab198d;
    ram_cell[     730] = 32'h1e8989ac;
    ram_cell[     731] = 32'h3f5846a3;
    ram_cell[     732] = 32'h39440f2e;
    ram_cell[     733] = 32'h29c8d58f;
    ram_cell[     734] = 32'h896b5e36;
    ram_cell[     735] = 32'h66b5f21b;
    ram_cell[     736] = 32'h0a7c9566;
    ram_cell[     737] = 32'h8a09b43c;
    ram_cell[     738] = 32'h9aad9dd9;
    ram_cell[     739] = 32'h7daac118;
    ram_cell[     740] = 32'h269a816b;
    ram_cell[     741] = 32'h1b9c4d64;
    ram_cell[     742] = 32'h8f2174b8;
    ram_cell[     743] = 32'h60bec763;
    ram_cell[     744] = 32'h23974052;
    ram_cell[     745] = 32'h4b67908a;
    ram_cell[     746] = 32'h05c49c4b;
    ram_cell[     747] = 32'ha9cba522;
    ram_cell[     748] = 32'hd30e6c9f;
    ram_cell[     749] = 32'h54e4c631;
    ram_cell[     750] = 32'h85a6f7c5;
    ram_cell[     751] = 32'h64891ba2;
    ram_cell[     752] = 32'he2245ecc;
    ram_cell[     753] = 32'h8a898096;
    ram_cell[     754] = 32'h0604354a;
    ram_cell[     755] = 32'h634f02ef;
    ram_cell[     756] = 32'hbecfa615;
    ram_cell[     757] = 32'h28ba327c;
    ram_cell[     758] = 32'h654ea693;
    ram_cell[     759] = 32'h34da2a3b;
    ram_cell[     760] = 32'hfa7a6ff7;
    ram_cell[     761] = 32'h7e289ea3;
    ram_cell[     762] = 32'h66129b63;
    ram_cell[     763] = 32'h6859e6cb;
    ram_cell[     764] = 32'h441a5ea7;
    ram_cell[     765] = 32'h4ce3092b;
    ram_cell[     766] = 32'h41840a9e;
    ram_cell[     767] = 32'h48a53fa0;
end

endmodule

