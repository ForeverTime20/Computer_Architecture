
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h3d34fd39;
    ram_cell[       1] = 32'h0;  // 32'hadce6b84;
    ram_cell[       2] = 32'h0;  // 32'h9ad0a6d3;
    ram_cell[       3] = 32'h0;  // 32'h4e59d51a;
    ram_cell[       4] = 32'h0;  // 32'h8804bf86;
    ram_cell[       5] = 32'h0;  // 32'hb1108b82;
    ram_cell[       6] = 32'h0;  // 32'hf99de8d0;
    ram_cell[       7] = 32'h0;  // 32'hf0bda0ef;
    ram_cell[       8] = 32'h0;  // 32'hba151d9d;
    ram_cell[       9] = 32'h0;  // 32'h568d438c;
    ram_cell[      10] = 32'h0;  // 32'hb56c3d37;
    ram_cell[      11] = 32'h0;  // 32'h5a4cb756;
    ram_cell[      12] = 32'h0;  // 32'heb78c1d5;
    ram_cell[      13] = 32'h0;  // 32'h7c9ca67e;
    ram_cell[      14] = 32'h0;  // 32'h7dd4b0de;
    ram_cell[      15] = 32'h0;  // 32'h85a0971c;
    ram_cell[      16] = 32'h0;  // 32'hf847401c;
    ram_cell[      17] = 32'h0;  // 32'h14d89913;
    ram_cell[      18] = 32'h0;  // 32'h279cdee8;
    ram_cell[      19] = 32'h0;  // 32'hb7dd0f8e;
    ram_cell[      20] = 32'h0;  // 32'heba5c9a0;
    ram_cell[      21] = 32'h0;  // 32'h81be77e2;
    ram_cell[      22] = 32'h0;  // 32'h9e13bc62;
    ram_cell[      23] = 32'h0;  // 32'hed7a227e;
    ram_cell[      24] = 32'h0;  // 32'h6ed25be1;
    ram_cell[      25] = 32'h0;  // 32'hfe374f5d;
    ram_cell[      26] = 32'h0;  // 32'h246e05ce;
    ram_cell[      27] = 32'h0;  // 32'hc81dee6c;
    ram_cell[      28] = 32'h0;  // 32'ha24c8ea3;
    ram_cell[      29] = 32'h0;  // 32'h19af0b9f;
    ram_cell[      30] = 32'h0;  // 32'h558ace7c;
    ram_cell[      31] = 32'h0;  // 32'h93810b98;
    ram_cell[      32] = 32'h0;  // 32'h8463be25;
    ram_cell[      33] = 32'h0;  // 32'hba2802ef;
    ram_cell[      34] = 32'h0;  // 32'hafe89893;
    ram_cell[      35] = 32'h0;  // 32'h5b422ec1;
    ram_cell[      36] = 32'h0;  // 32'hd5c327f1;
    ram_cell[      37] = 32'h0;  // 32'hab739b5e;
    ram_cell[      38] = 32'h0;  // 32'h39628eea;
    ram_cell[      39] = 32'h0;  // 32'hf9cdcfac;
    ram_cell[      40] = 32'h0;  // 32'h7cb1e321;
    ram_cell[      41] = 32'h0;  // 32'h90505b03;
    ram_cell[      42] = 32'h0;  // 32'hcc5e7808;
    ram_cell[      43] = 32'h0;  // 32'h884c7228;
    ram_cell[      44] = 32'h0;  // 32'h72d1fb92;
    ram_cell[      45] = 32'h0;  // 32'h3925f635;
    ram_cell[      46] = 32'h0;  // 32'ha4febd9c;
    ram_cell[      47] = 32'h0;  // 32'h8f0e0c1c;
    ram_cell[      48] = 32'h0;  // 32'h6ad0a82c;
    ram_cell[      49] = 32'h0;  // 32'hb78ab1bf;
    ram_cell[      50] = 32'h0;  // 32'h0427a70f;
    ram_cell[      51] = 32'h0;  // 32'hb1cf274f;
    ram_cell[      52] = 32'h0;  // 32'he6a3964c;
    ram_cell[      53] = 32'h0;  // 32'h3ee8b5ce;
    ram_cell[      54] = 32'h0;  // 32'h87a06727;
    ram_cell[      55] = 32'h0;  // 32'h16f9a70e;
    ram_cell[      56] = 32'h0;  // 32'h2ac84d16;
    ram_cell[      57] = 32'h0;  // 32'hc405b6de;
    ram_cell[      58] = 32'h0;  // 32'he6219dd8;
    ram_cell[      59] = 32'h0;  // 32'ha4e42d6e;
    ram_cell[      60] = 32'h0;  // 32'h24e47248;
    ram_cell[      61] = 32'h0;  // 32'ha6d092e8;
    ram_cell[      62] = 32'h0;  // 32'hb5d62b56;
    ram_cell[      63] = 32'h0;  // 32'hce9bb880;
    ram_cell[      64] = 32'h0;  // 32'h30db21f5;
    ram_cell[      65] = 32'h0;  // 32'hc7e7f787;
    ram_cell[      66] = 32'h0;  // 32'hf580d362;
    ram_cell[      67] = 32'h0;  // 32'h804fbe22;
    ram_cell[      68] = 32'h0;  // 32'h3e036c9a;
    ram_cell[      69] = 32'h0;  // 32'h71b0d341;
    ram_cell[      70] = 32'h0;  // 32'h4ea45bf1;
    ram_cell[      71] = 32'h0;  // 32'h9e674c15;
    ram_cell[      72] = 32'h0;  // 32'h8f40c6e7;
    ram_cell[      73] = 32'h0;  // 32'h2ff17c5d;
    ram_cell[      74] = 32'h0;  // 32'h6d356ebb;
    ram_cell[      75] = 32'h0;  // 32'h56eed951;
    ram_cell[      76] = 32'h0;  // 32'hac649740;
    ram_cell[      77] = 32'h0;  // 32'h2f5d9598;
    ram_cell[      78] = 32'h0;  // 32'hb2fa82c8;
    ram_cell[      79] = 32'h0;  // 32'hb51976d2;
    ram_cell[      80] = 32'h0;  // 32'h5bab9945;
    ram_cell[      81] = 32'h0;  // 32'h500fcd7a;
    ram_cell[      82] = 32'h0;  // 32'hde683644;
    ram_cell[      83] = 32'h0;  // 32'hdc0a4246;
    ram_cell[      84] = 32'h0;  // 32'hbc98f62a;
    ram_cell[      85] = 32'h0;  // 32'h4cc105e5;
    ram_cell[      86] = 32'h0;  // 32'h70a9ff32;
    ram_cell[      87] = 32'h0;  // 32'h229f29fa;
    ram_cell[      88] = 32'h0;  // 32'hb6ed6345;
    ram_cell[      89] = 32'h0;  // 32'h30640798;
    ram_cell[      90] = 32'h0;  // 32'h6c538358;
    ram_cell[      91] = 32'h0;  // 32'h9afc3fa4;
    ram_cell[      92] = 32'h0;  // 32'h959325ea;
    ram_cell[      93] = 32'h0;  // 32'hfabd78d4;
    ram_cell[      94] = 32'h0;  // 32'h6123a16c;
    ram_cell[      95] = 32'h0;  // 32'h5dc28110;
    ram_cell[      96] = 32'h0;  // 32'h6607e33f;
    ram_cell[      97] = 32'h0;  // 32'h43b9ffbe;
    ram_cell[      98] = 32'h0;  // 32'h73a569ad;
    ram_cell[      99] = 32'h0;  // 32'h33fe9470;
    ram_cell[     100] = 32'h0;  // 32'hb4ed70c6;
    ram_cell[     101] = 32'h0;  // 32'h3c7fb3e6;
    ram_cell[     102] = 32'h0;  // 32'he113abec;
    ram_cell[     103] = 32'h0;  // 32'had2cc481;
    ram_cell[     104] = 32'h0;  // 32'h256e850c;
    ram_cell[     105] = 32'h0;  // 32'h05ff06b1;
    ram_cell[     106] = 32'h0;  // 32'hbccbcea2;
    ram_cell[     107] = 32'h0;  // 32'hb025c848;
    ram_cell[     108] = 32'h0;  // 32'hc9d5aa52;
    ram_cell[     109] = 32'h0;  // 32'hfe0646f1;
    ram_cell[     110] = 32'h0;  // 32'he996f44d;
    ram_cell[     111] = 32'h0;  // 32'ha2fdd9f0;
    ram_cell[     112] = 32'h0;  // 32'hdbb40bbf;
    ram_cell[     113] = 32'h0;  // 32'h1900e5c9;
    ram_cell[     114] = 32'h0;  // 32'hf0e26819;
    ram_cell[     115] = 32'h0;  // 32'h74f56601;
    ram_cell[     116] = 32'h0;  // 32'h50b3ee6c;
    ram_cell[     117] = 32'h0;  // 32'h8783ae22;
    ram_cell[     118] = 32'h0;  // 32'hae6775d0;
    ram_cell[     119] = 32'h0;  // 32'hb94bd3c6;
    ram_cell[     120] = 32'h0;  // 32'haaeee287;
    ram_cell[     121] = 32'h0;  // 32'h8adda877;
    ram_cell[     122] = 32'h0;  // 32'h0b9e3a11;
    ram_cell[     123] = 32'h0;  // 32'h920e049e;
    ram_cell[     124] = 32'h0;  // 32'h4e614005;
    ram_cell[     125] = 32'h0;  // 32'h13288054;
    ram_cell[     126] = 32'h0;  // 32'h06caef88;
    ram_cell[     127] = 32'h0;  // 32'h3ca8375b;
    ram_cell[     128] = 32'h0;  // 32'h683cf034;
    ram_cell[     129] = 32'h0;  // 32'hde5debc1;
    ram_cell[     130] = 32'h0;  // 32'h579b9390;
    ram_cell[     131] = 32'h0;  // 32'h2982dba8;
    ram_cell[     132] = 32'h0;  // 32'h7278c9cd;
    ram_cell[     133] = 32'h0;  // 32'h5106cab1;
    ram_cell[     134] = 32'h0;  // 32'hfd07bf38;
    ram_cell[     135] = 32'h0;  // 32'h19ba1ff1;
    ram_cell[     136] = 32'h0;  // 32'hc32e81a1;
    ram_cell[     137] = 32'h0;  // 32'h7f6dad72;
    ram_cell[     138] = 32'h0;  // 32'hf2655918;
    ram_cell[     139] = 32'h0;  // 32'ha04fb8f9;
    ram_cell[     140] = 32'h0;  // 32'h07d86553;
    ram_cell[     141] = 32'h0;  // 32'hb5721a72;
    ram_cell[     142] = 32'h0;  // 32'hd8237a6b;
    ram_cell[     143] = 32'h0;  // 32'h6b57e418;
    ram_cell[     144] = 32'h0;  // 32'heecbf30c;
    ram_cell[     145] = 32'h0;  // 32'hf9b2ca60;
    ram_cell[     146] = 32'h0;  // 32'h836b7176;
    ram_cell[     147] = 32'h0;  // 32'h07f84c38;
    ram_cell[     148] = 32'h0;  // 32'hf719be9c;
    ram_cell[     149] = 32'h0;  // 32'h58459056;
    ram_cell[     150] = 32'h0;  // 32'he4b94c9e;
    ram_cell[     151] = 32'h0;  // 32'h77650453;
    ram_cell[     152] = 32'h0;  // 32'hcc129c27;
    ram_cell[     153] = 32'h0;  // 32'h96bb1c00;
    ram_cell[     154] = 32'h0;  // 32'h82719d1a;
    ram_cell[     155] = 32'h0;  // 32'h20f4505e;
    ram_cell[     156] = 32'h0;  // 32'h5b96953c;
    ram_cell[     157] = 32'h0;  // 32'h7dd12b95;
    ram_cell[     158] = 32'h0;  // 32'h4e21dbf1;
    ram_cell[     159] = 32'h0;  // 32'h1c873955;
    ram_cell[     160] = 32'h0;  // 32'ha5ddf14e;
    ram_cell[     161] = 32'h0;  // 32'hc4d31c3a;
    ram_cell[     162] = 32'h0;  // 32'h50cd1ad2;
    ram_cell[     163] = 32'h0;  // 32'h1cd90368;
    ram_cell[     164] = 32'h0;  // 32'hc3918f48;
    ram_cell[     165] = 32'h0;  // 32'h5766af64;
    ram_cell[     166] = 32'h0;  // 32'h479b0833;
    ram_cell[     167] = 32'h0;  // 32'h761a0114;
    ram_cell[     168] = 32'h0;  // 32'h63152327;
    ram_cell[     169] = 32'h0;  // 32'hdf42fd8e;
    ram_cell[     170] = 32'h0;  // 32'hb20cf7f3;
    ram_cell[     171] = 32'h0;  // 32'h7b42a947;
    ram_cell[     172] = 32'h0;  // 32'h25eafa12;
    ram_cell[     173] = 32'h0;  // 32'hb6e639ce;
    ram_cell[     174] = 32'h0;  // 32'h41c509c5;
    ram_cell[     175] = 32'h0;  // 32'h27b6c2f9;
    ram_cell[     176] = 32'h0;  // 32'hb638fa7b;
    ram_cell[     177] = 32'h0;  // 32'hb33c9b94;
    ram_cell[     178] = 32'h0;  // 32'ha3c58a30;
    ram_cell[     179] = 32'h0;  // 32'h420d4c38;
    ram_cell[     180] = 32'h0;  // 32'hc0ccbeac;
    ram_cell[     181] = 32'h0;  // 32'h1cd44375;
    ram_cell[     182] = 32'h0;  // 32'hc118c721;
    ram_cell[     183] = 32'h0;  // 32'h7f864e78;
    ram_cell[     184] = 32'h0;  // 32'h5f1c2cfe;
    ram_cell[     185] = 32'h0;  // 32'hd9aedbcf;
    ram_cell[     186] = 32'h0;  // 32'h8d575e0a;
    ram_cell[     187] = 32'h0;  // 32'hbd95a4e7;
    ram_cell[     188] = 32'h0;  // 32'hc2dd84e2;
    ram_cell[     189] = 32'h0;  // 32'hdf762a93;
    ram_cell[     190] = 32'h0;  // 32'h3e1d675d;
    ram_cell[     191] = 32'h0;  // 32'hbb41d064;
    ram_cell[     192] = 32'h0;  // 32'h36153d6e;
    ram_cell[     193] = 32'h0;  // 32'h5d6f613f;
    ram_cell[     194] = 32'h0;  // 32'h837a0c71;
    ram_cell[     195] = 32'h0;  // 32'h3c4ff6a3;
    ram_cell[     196] = 32'h0;  // 32'h94bdfcae;
    ram_cell[     197] = 32'h0;  // 32'h6a05969c;
    ram_cell[     198] = 32'h0;  // 32'h1cfe1d47;
    ram_cell[     199] = 32'h0;  // 32'h49e28178;
    ram_cell[     200] = 32'h0;  // 32'h8b18f5b2;
    ram_cell[     201] = 32'h0;  // 32'h38044ca7;
    ram_cell[     202] = 32'h0;  // 32'h6837c925;
    ram_cell[     203] = 32'h0;  // 32'h4c263562;
    ram_cell[     204] = 32'h0;  // 32'h52514ac1;
    ram_cell[     205] = 32'h0;  // 32'h6055a1e9;
    ram_cell[     206] = 32'h0;  // 32'h7e71cb06;
    ram_cell[     207] = 32'h0;  // 32'h2924bf05;
    ram_cell[     208] = 32'h0;  // 32'ha88f5262;
    ram_cell[     209] = 32'h0;  // 32'he6068408;
    ram_cell[     210] = 32'h0;  // 32'h24d2644c;
    ram_cell[     211] = 32'h0;  // 32'hee890cb7;
    ram_cell[     212] = 32'h0;  // 32'hc480bcb3;
    ram_cell[     213] = 32'h0;  // 32'hdd310f52;
    ram_cell[     214] = 32'h0;  // 32'h56512759;
    ram_cell[     215] = 32'h0;  // 32'h0c936365;
    ram_cell[     216] = 32'h0;  // 32'h7aa30c9b;
    ram_cell[     217] = 32'h0;  // 32'h45184363;
    ram_cell[     218] = 32'h0;  // 32'h1c2eefea;
    ram_cell[     219] = 32'h0;  // 32'hed083ce4;
    ram_cell[     220] = 32'h0;  // 32'ha8f2e5e8;
    ram_cell[     221] = 32'h0;  // 32'hf33bfc71;
    ram_cell[     222] = 32'h0;  // 32'h2b20b170;
    ram_cell[     223] = 32'h0;  // 32'he4da7074;
    ram_cell[     224] = 32'h0;  // 32'h4d56da2a;
    ram_cell[     225] = 32'h0;  // 32'h3144c547;
    ram_cell[     226] = 32'h0;  // 32'h7bb382bf;
    ram_cell[     227] = 32'h0;  // 32'hea0e970d;
    ram_cell[     228] = 32'h0;  // 32'hd7cb168d;
    ram_cell[     229] = 32'h0;  // 32'h8b2fdfd1;
    ram_cell[     230] = 32'h0;  // 32'h4617445f;
    ram_cell[     231] = 32'h0;  // 32'hb9802a78;
    ram_cell[     232] = 32'h0;  // 32'h979c2437;
    ram_cell[     233] = 32'h0;  // 32'hae96a44f;
    ram_cell[     234] = 32'h0;  // 32'h333fd7f9;
    ram_cell[     235] = 32'h0;  // 32'hbd4d51e0;
    ram_cell[     236] = 32'h0;  // 32'h4db873b8;
    ram_cell[     237] = 32'h0;  // 32'hb5550b48;
    ram_cell[     238] = 32'h0;  // 32'hce3590ce;
    ram_cell[     239] = 32'h0;  // 32'hb7adca6e;
    ram_cell[     240] = 32'h0;  // 32'hd395b716;
    ram_cell[     241] = 32'h0;  // 32'hf3647f8c;
    ram_cell[     242] = 32'h0;  // 32'h427c8517;
    ram_cell[     243] = 32'h0;  // 32'h96e96027;
    ram_cell[     244] = 32'h0;  // 32'hf7344cad;
    ram_cell[     245] = 32'h0;  // 32'h3e3eeca6;
    ram_cell[     246] = 32'h0;  // 32'h896367f9;
    ram_cell[     247] = 32'h0;  // 32'hc91c9df5;
    ram_cell[     248] = 32'h0;  // 32'ha416f473;
    ram_cell[     249] = 32'h0;  // 32'h8add508c;
    ram_cell[     250] = 32'h0;  // 32'h7a488b4d;
    ram_cell[     251] = 32'h0;  // 32'hd9ecc0aa;
    ram_cell[     252] = 32'h0;  // 32'h60833406;
    ram_cell[     253] = 32'h0;  // 32'h38004a5a;
    ram_cell[     254] = 32'h0;  // 32'h9d1684e7;
    ram_cell[     255] = 32'h0;  // 32'h00c29064;
    // src matrix A
    ram_cell[     256] = 32'ha3cd3575;
    ram_cell[     257] = 32'h39ab396f;
    ram_cell[     258] = 32'h5d79c425;
    ram_cell[     259] = 32'he21ff36a;
    ram_cell[     260] = 32'hb58fa9ea;
    ram_cell[     261] = 32'h76ab2a86;
    ram_cell[     262] = 32'h92e3d264;
    ram_cell[     263] = 32'h2e4b30a5;
    ram_cell[     264] = 32'hafd7f8c2;
    ram_cell[     265] = 32'he7f4a594;
    ram_cell[     266] = 32'h4993d6f5;
    ram_cell[     267] = 32'h991b4668;
    ram_cell[     268] = 32'haacf3fe9;
    ram_cell[     269] = 32'h1bc585b7;
    ram_cell[     270] = 32'h0345a3da;
    ram_cell[     271] = 32'h5d18be9f;
    ram_cell[     272] = 32'hcdf45e91;
    ram_cell[     273] = 32'h50a43a1e;
    ram_cell[     274] = 32'h00b36417;
    ram_cell[     275] = 32'h67a48115;
    ram_cell[     276] = 32'heedaf701;
    ram_cell[     277] = 32'h707fddee;
    ram_cell[     278] = 32'h82ae0170;
    ram_cell[     279] = 32'hbbf3d41a;
    ram_cell[     280] = 32'h4b19b987;
    ram_cell[     281] = 32'h320c2649;
    ram_cell[     282] = 32'h54702032;
    ram_cell[     283] = 32'h0b9b3f38;
    ram_cell[     284] = 32'h4f5bcff2;
    ram_cell[     285] = 32'hb7908c79;
    ram_cell[     286] = 32'hf8765135;
    ram_cell[     287] = 32'hfd2d4dec;
    ram_cell[     288] = 32'h06db2a8a;
    ram_cell[     289] = 32'h1d685101;
    ram_cell[     290] = 32'h16026470;
    ram_cell[     291] = 32'hdd9d20c4;
    ram_cell[     292] = 32'hc6005aa6;
    ram_cell[     293] = 32'hd9ee5aac;
    ram_cell[     294] = 32'h53c416e1;
    ram_cell[     295] = 32'h996586d5;
    ram_cell[     296] = 32'hac53b25c;
    ram_cell[     297] = 32'hf215ba50;
    ram_cell[     298] = 32'hdbdd99a7;
    ram_cell[     299] = 32'h2e327f9b;
    ram_cell[     300] = 32'hca46787d;
    ram_cell[     301] = 32'h7c12e037;
    ram_cell[     302] = 32'h8ef090b0;
    ram_cell[     303] = 32'h13873d96;
    ram_cell[     304] = 32'hf82d0336;
    ram_cell[     305] = 32'h42d46df1;
    ram_cell[     306] = 32'heb40946b;
    ram_cell[     307] = 32'h7012eb26;
    ram_cell[     308] = 32'ha89a2854;
    ram_cell[     309] = 32'hd1760369;
    ram_cell[     310] = 32'h460781f3;
    ram_cell[     311] = 32'h7952583d;
    ram_cell[     312] = 32'h4e1b3eb9;
    ram_cell[     313] = 32'hcc3f93c8;
    ram_cell[     314] = 32'h19603990;
    ram_cell[     315] = 32'hd714e726;
    ram_cell[     316] = 32'hd9f61ce7;
    ram_cell[     317] = 32'h2a7b9b08;
    ram_cell[     318] = 32'h0fb39409;
    ram_cell[     319] = 32'ha7f394b8;
    ram_cell[     320] = 32'he881e52e;
    ram_cell[     321] = 32'hb3c5b6e0;
    ram_cell[     322] = 32'he04bbafa;
    ram_cell[     323] = 32'hdd5c185e;
    ram_cell[     324] = 32'h52d78160;
    ram_cell[     325] = 32'hbe471f96;
    ram_cell[     326] = 32'h74253642;
    ram_cell[     327] = 32'hc771781f;
    ram_cell[     328] = 32'h37cb6b78;
    ram_cell[     329] = 32'h18a5feb2;
    ram_cell[     330] = 32'h2f669462;
    ram_cell[     331] = 32'h47ab1d8b;
    ram_cell[     332] = 32'haa8d691e;
    ram_cell[     333] = 32'he5f11978;
    ram_cell[     334] = 32'h51f3a71c;
    ram_cell[     335] = 32'h07b0ed13;
    ram_cell[     336] = 32'hd0b7e868;
    ram_cell[     337] = 32'h4234f3b9;
    ram_cell[     338] = 32'hdcf98ef4;
    ram_cell[     339] = 32'h9acc965b;
    ram_cell[     340] = 32'h3c67dfff;
    ram_cell[     341] = 32'h1eddad6e;
    ram_cell[     342] = 32'h93328e1b;
    ram_cell[     343] = 32'ha43ee105;
    ram_cell[     344] = 32'h69e25e35;
    ram_cell[     345] = 32'h4b288568;
    ram_cell[     346] = 32'h93548c83;
    ram_cell[     347] = 32'h4d589428;
    ram_cell[     348] = 32'hf120344b;
    ram_cell[     349] = 32'habfd765a;
    ram_cell[     350] = 32'h05b8a68e;
    ram_cell[     351] = 32'h4065d591;
    ram_cell[     352] = 32'h7f137d2c;
    ram_cell[     353] = 32'hf40af52f;
    ram_cell[     354] = 32'hf3672ca9;
    ram_cell[     355] = 32'h522e205c;
    ram_cell[     356] = 32'h2769503a;
    ram_cell[     357] = 32'had7e1a44;
    ram_cell[     358] = 32'h0551966f;
    ram_cell[     359] = 32'h991e5b9f;
    ram_cell[     360] = 32'hd82d8b61;
    ram_cell[     361] = 32'h10d949e8;
    ram_cell[     362] = 32'hc1c8f950;
    ram_cell[     363] = 32'h36e4cb04;
    ram_cell[     364] = 32'h4c6123a4;
    ram_cell[     365] = 32'he17b853f;
    ram_cell[     366] = 32'h5e120e82;
    ram_cell[     367] = 32'h6687c584;
    ram_cell[     368] = 32'h95c10b0d;
    ram_cell[     369] = 32'hae5eb768;
    ram_cell[     370] = 32'h9e35fd32;
    ram_cell[     371] = 32'h6421cbcd;
    ram_cell[     372] = 32'h47df016f;
    ram_cell[     373] = 32'hb2a2fa15;
    ram_cell[     374] = 32'ha176c616;
    ram_cell[     375] = 32'h4c178ab1;
    ram_cell[     376] = 32'h35759bce;
    ram_cell[     377] = 32'h02a0bad6;
    ram_cell[     378] = 32'h42901bba;
    ram_cell[     379] = 32'h772d507c;
    ram_cell[     380] = 32'hec14d0ef;
    ram_cell[     381] = 32'hec20ee3a;
    ram_cell[     382] = 32'h331387b9;
    ram_cell[     383] = 32'h4fe92039;
    ram_cell[     384] = 32'h3c94d474;
    ram_cell[     385] = 32'hfdd64e95;
    ram_cell[     386] = 32'h3054d76e;
    ram_cell[     387] = 32'hee378e1b;
    ram_cell[     388] = 32'h163aff12;
    ram_cell[     389] = 32'he55b30bf;
    ram_cell[     390] = 32'h62ce0f05;
    ram_cell[     391] = 32'h14db444e;
    ram_cell[     392] = 32'h84f0d8fe;
    ram_cell[     393] = 32'h379feafa;
    ram_cell[     394] = 32'h45da4de0;
    ram_cell[     395] = 32'h17a817fb;
    ram_cell[     396] = 32'h5966b0aa;
    ram_cell[     397] = 32'h27aa9f58;
    ram_cell[     398] = 32'h0dc85fdc;
    ram_cell[     399] = 32'h44d0d8ac;
    ram_cell[     400] = 32'h110647be;
    ram_cell[     401] = 32'h820a3472;
    ram_cell[     402] = 32'hb49f5819;
    ram_cell[     403] = 32'hd6fddc47;
    ram_cell[     404] = 32'hff154594;
    ram_cell[     405] = 32'h2916a565;
    ram_cell[     406] = 32'hb0f4526c;
    ram_cell[     407] = 32'hec9b535c;
    ram_cell[     408] = 32'h480eae2e;
    ram_cell[     409] = 32'hd80260d8;
    ram_cell[     410] = 32'hb3be2937;
    ram_cell[     411] = 32'h8414a355;
    ram_cell[     412] = 32'hbfe0298e;
    ram_cell[     413] = 32'h4a1c758c;
    ram_cell[     414] = 32'h0462c5f3;
    ram_cell[     415] = 32'hed2b87be;
    ram_cell[     416] = 32'hf165e288;
    ram_cell[     417] = 32'h6889a0d1;
    ram_cell[     418] = 32'h7ce0d84d;
    ram_cell[     419] = 32'h75ab1b8f;
    ram_cell[     420] = 32'h9d28d2d7;
    ram_cell[     421] = 32'h40113d4a;
    ram_cell[     422] = 32'h94950126;
    ram_cell[     423] = 32'h8b3ab1e7;
    ram_cell[     424] = 32'hdb6e4027;
    ram_cell[     425] = 32'hbc884a3b;
    ram_cell[     426] = 32'h8ca31f62;
    ram_cell[     427] = 32'hb6737208;
    ram_cell[     428] = 32'hd7671055;
    ram_cell[     429] = 32'hed0fbff1;
    ram_cell[     430] = 32'hda8da4b6;
    ram_cell[     431] = 32'h00443785;
    ram_cell[     432] = 32'hacacc14c;
    ram_cell[     433] = 32'h7e924e01;
    ram_cell[     434] = 32'h9fbe70f3;
    ram_cell[     435] = 32'h24e88720;
    ram_cell[     436] = 32'heb1d1447;
    ram_cell[     437] = 32'h7eba1988;
    ram_cell[     438] = 32'h0d31295f;
    ram_cell[     439] = 32'he2bce333;
    ram_cell[     440] = 32'h178397d1;
    ram_cell[     441] = 32'h681772c6;
    ram_cell[     442] = 32'h2147cfc4;
    ram_cell[     443] = 32'h47433006;
    ram_cell[     444] = 32'h76853886;
    ram_cell[     445] = 32'h66bd0886;
    ram_cell[     446] = 32'h3437ab54;
    ram_cell[     447] = 32'h5638902f;
    ram_cell[     448] = 32'hb0b30741;
    ram_cell[     449] = 32'ha23b8be0;
    ram_cell[     450] = 32'h3fbde09a;
    ram_cell[     451] = 32'h01800c3a;
    ram_cell[     452] = 32'hc76ebee5;
    ram_cell[     453] = 32'hb297393f;
    ram_cell[     454] = 32'h920d600e;
    ram_cell[     455] = 32'hdfab1e92;
    ram_cell[     456] = 32'h695aaaff;
    ram_cell[     457] = 32'hda627e4e;
    ram_cell[     458] = 32'haca3e832;
    ram_cell[     459] = 32'hfdc9bdf4;
    ram_cell[     460] = 32'hde93f26f;
    ram_cell[     461] = 32'h4b619dd8;
    ram_cell[     462] = 32'h3ab347ee;
    ram_cell[     463] = 32'h2813cf3e;
    ram_cell[     464] = 32'h6afef99a;
    ram_cell[     465] = 32'h50bea73b;
    ram_cell[     466] = 32'h8313a916;
    ram_cell[     467] = 32'h60b9486d;
    ram_cell[     468] = 32'hd46ccc3e;
    ram_cell[     469] = 32'h32c7adc9;
    ram_cell[     470] = 32'h88185f7f;
    ram_cell[     471] = 32'hf1ac7d43;
    ram_cell[     472] = 32'ha7f3f0d5;
    ram_cell[     473] = 32'hdc851389;
    ram_cell[     474] = 32'h0c80132d;
    ram_cell[     475] = 32'h14048bb8;
    ram_cell[     476] = 32'hd616460d;
    ram_cell[     477] = 32'hf3580232;
    ram_cell[     478] = 32'h55db1d51;
    ram_cell[     479] = 32'ha4eba88c;
    ram_cell[     480] = 32'hff2e14a6;
    ram_cell[     481] = 32'h0f9ab187;
    ram_cell[     482] = 32'h85b1d19b;
    ram_cell[     483] = 32'h1374ba2a;
    ram_cell[     484] = 32'h715745c6;
    ram_cell[     485] = 32'h5dd08619;
    ram_cell[     486] = 32'h71722b07;
    ram_cell[     487] = 32'hea8c4857;
    ram_cell[     488] = 32'ha8f7ccdb;
    ram_cell[     489] = 32'hf9ee643c;
    ram_cell[     490] = 32'h169f46e9;
    ram_cell[     491] = 32'ha3f71348;
    ram_cell[     492] = 32'hcbad68d7;
    ram_cell[     493] = 32'h806172f0;
    ram_cell[     494] = 32'hb1171b22;
    ram_cell[     495] = 32'h0d5c22b5;
    ram_cell[     496] = 32'haf84e8e7;
    ram_cell[     497] = 32'h1d4e5bbe;
    ram_cell[     498] = 32'h8a5035e5;
    ram_cell[     499] = 32'h288d4bdd;
    ram_cell[     500] = 32'h0f32d207;
    ram_cell[     501] = 32'hcef331fb;
    ram_cell[     502] = 32'h377e2bc7;
    ram_cell[     503] = 32'h76aa60f2;
    ram_cell[     504] = 32'h585a4044;
    ram_cell[     505] = 32'hcf47af36;
    ram_cell[     506] = 32'h9f29bcb5;
    ram_cell[     507] = 32'hd2748abb;
    ram_cell[     508] = 32'h1fc22e73;
    ram_cell[     509] = 32'h9973eae0;
    ram_cell[     510] = 32'he2e95607;
    ram_cell[     511] = 32'h27df63f8;
    // src matrix B
    ram_cell[     512] = 32'h119e988d;
    ram_cell[     513] = 32'h8a4f2c45;
    ram_cell[     514] = 32'h042eb84f;
    ram_cell[     515] = 32'h0fc146d5;
    ram_cell[     516] = 32'h832e86bc;
    ram_cell[     517] = 32'h0375129f;
    ram_cell[     518] = 32'h7746e004;
    ram_cell[     519] = 32'h66265eaa;
    ram_cell[     520] = 32'h1ea56d57;
    ram_cell[     521] = 32'h4a276280;
    ram_cell[     522] = 32'hb45709f9;
    ram_cell[     523] = 32'h9227480e;
    ram_cell[     524] = 32'h2efea336;
    ram_cell[     525] = 32'h6be1f239;
    ram_cell[     526] = 32'h6aa1b6f4;
    ram_cell[     527] = 32'he4cc6628;
    ram_cell[     528] = 32'h153e2fba;
    ram_cell[     529] = 32'h2bec5d1d;
    ram_cell[     530] = 32'h75f80c38;
    ram_cell[     531] = 32'h82a73d5f;
    ram_cell[     532] = 32'h554d3dcb;
    ram_cell[     533] = 32'hc6ccc007;
    ram_cell[     534] = 32'h93252d0d;
    ram_cell[     535] = 32'ha8ea4f1c;
    ram_cell[     536] = 32'ha7c0f9b5;
    ram_cell[     537] = 32'h535d3088;
    ram_cell[     538] = 32'had64dc9c;
    ram_cell[     539] = 32'h368c0dc4;
    ram_cell[     540] = 32'h3448faf8;
    ram_cell[     541] = 32'hc32a1d2d;
    ram_cell[     542] = 32'haf4e42d9;
    ram_cell[     543] = 32'hba4ce38c;
    ram_cell[     544] = 32'h4ae06d88;
    ram_cell[     545] = 32'ha7dbc8c4;
    ram_cell[     546] = 32'ha4739e80;
    ram_cell[     547] = 32'ha7f36155;
    ram_cell[     548] = 32'hd0bd7758;
    ram_cell[     549] = 32'h9c2e5343;
    ram_cell[     550] = 32'h0300d1d5;
    ram_cell[     551] = 32'h4573fe60;
    ram_cell[     552] = 32'hc94e8262;
    ram_cell[     553] = 32'h81230c57;
    ram_cell[     554] = 32'h347b621f;
    ram_cell[     555] = 32'h433c9e5f;
    ram_cell[     556] = 32'h1adee3c4;
    ram_cell[     557] = 32'h5a82f9be;
    ram_cell[     558] = 32'hae62dec4;
    ram_cell[     559] = 32'h4ca53316;
    ram_cell[     560] = 32'h9d75fcae;
    ram_cell[     561] = 32'h0a54b59a;
    ram_cell[     562] = 32'h799f9898;
    ram_cell[     563] = 32'h5853615d;
    ram_cell[     564] = 32'h05f5e63f;
    ram_cell[     565] = 32'h9a6c1587;
    ram_cell[     566] = 32'h6a3d4319;
    ram_cell[     567] = 32'h28d7cd24;
    ram_cell[     568] = 32'h0b3a6295;
    ram_cell[     569] = 32'h3e45db78;
    ram_cell[     570] = 32'h2bb36867;
    ram_cell[     571] = 32'h23395f4b;
    ram_cell[     572] = 32'h8802c875;
    ram_cell[     573] = 32'h86adf0cc;
    ram_cell[     574] = 32'hccf99965;
    ram_cell[     575] = 32'h6354abe1;
    ram_cell[     576] = 32'h2de1f139;
    ram_cell[     577] = 32'h3bc92f15;
    ram_cell[     578] = 32'hc36f19fc;
    ram_cell[     579] = 32'h96852019;
    ram_cell[     580] = 32'h30cfa563;
    ram_cell[     581] = 32'h98d55d6f;
    ram_cell[     582] = 32'h75605e4b;
    ram_cell[     583] = 32'h8eb410ae;
    ram_cell[     584] = 32'ha777d7a0;
    ram_cell[     585] = 32'h69d82b39;
    ram_cell[     586] = 32'h7902f7ba;
    ram_cell[     587] = 32'hf7e1e4f1;
    ram_cell[     588] = 32'hba398912;
    ram_cell[     589] = 32'h3412fb51;
    ram_cell[     590] = 32'h561cffa7;
    ram_cell[     591] = 32'hb480ca23;
    ram_cell[     592] = 32'hf42eb3bc;
    ram_cell[     593] = 32'h81ea94f4;
    ram_cell[     594] = 32'h550cd871;
    ram_cell[     595] = 32'hbbeaee5c;
    ram_cell[     596] = 32'h4e8304f7;
    ram_cell[     597] = 32'h8b84bc3d;
    ram_cell[     598] = 32'h00736206;
    ram_cell[     599] = 32'h10855118;
    ram_cell[     600] = 32'h8a8a04fd;
    ram_cell[     601] = 32'h0266a96d;
    ram_cell[     602] = 32'h32045099;
    ram_cell[     603] = 32'h63c75c1b;
    ram_cell[     604] = 32'h9bd4b1c3;
    ram_cell[     605] = 32'h2c804dd5;
    ram_cell[     606] = 32'hd3408608;
    ram_cell[     607] = 32'hc3b91bc0;
    ram_cell[     608] = 32'hf59e2e6f;
    ram_cell[     609] = 32'h2e86e1ce;
    ram_cell[     610] = 32'hb9fcfe8c;
    ram_cell[     611] = 32'haba6afc5;
    ram_cell[     612] = 32'h76441ba8;
    ram_cell[     613] = 32'hcd2eb2a6;
    ram_cell[     614] = 32'h3d3c34a7;
    ram_cell[     615] = 32'h5659209a;
    ram_cell[     616] = 32'h9c3dd759;
    ram_cell[     617] = 32'h4bd6e8e9;
    ram_cell[     618] = 32'he2362bef;
    ram_cell[     619] = 32'hd2d3d940;
    ram_cell[     620] = 32'h42d570ab;
    ram_cell[     621] = 32'he0a71d16;
    ram_cell[     622] = 32'h57862966;
    ram_cell[     623] = 32'head1dbd0;
    ram_cell[     624] = 32'hbb46f3a7;
    ram_cell[     625] = 32'h34a902b3;
    ram_cell[     626] = 32'hbbfe5265;
    ram_cell[     627] = 32'hb71afab0;
    ram_cell[     628] = 32'hc4bcce5d;
    ram_cell[     629] = 32'h6943ff8f;
    ram_cell[     630] = 32'ha4017ead;
    ram_cell[     631] = 32'hef5527b6;
    ram_cell[     632] = 32'h9c33fcd7;
    ram_cell[     633] = 32'h0fe18b6c;
    ram_cell[     634] = 32'h9a12ba09;
    ram_cell[     635] = 32'hbad1db32;
    ram_cell[     636] = 32'h05974a8e;
    ram_cell[     637] = 32'hf4c57804;
    ram_cell[     638] = 32'h617585e6;
    ram_cell[     639] = 32'hf3205f56;
    ram_cell[     640] = 32'hc2735681;
    ram_cell[     641] = 32'h39a1c3a5;
    ram_cell[     642] = 32'h990159a5;
    ram_cell[     643] = 32'ha6199bd5;
    ram_cell[     644] = 32'h8914a36a;
    ram_cell[     645] = 32'hb2be0c27;
    ram_cell[     646] = 32'h60c2db5d;
    ram_cell[     647] = 32'h5df700de;
    ram_cell[     648] = 32'hc2a92584;
    ram_cell[     649] = 32'h0a705c1f;
    ram_cell[     650] = 32'h3660c2c8;
    ram_cell[     651] = 32'h42fd20bb;
    ram_cell[     652] = 32'h0f0c54ff;
    ram_cell[     653] = 32'h1f432497;
    ram_cell[     654] = 32'h28935ec0;
    ram_cell[     655] = 32'hc836ea44;
    ram_cell[     656] = 32'hf2a8abd7;
    ram_cell[     657] = 32'h002f28e9;
    ram_cell[     658] = 32'h9ecda88d;
    ram_cell[     659] = 32'h3a5e1896;
    ram_cell[     660] = 32'h23860d65;
    ram_cell[     661] = 32'h726ed0b4;
    ram_cell[     662] = 32'h433942be;
    ram_cell[     663] = 32'h7dbd5531;
    ram_cell[     664] = 32'h4b65233e;
    ram_cell[     665] = 32'h6566c11c;
    ram_cell[     666] = 32'h6ff677fb;
    ram_cell[     667] = 32'hbeb329b0;
    ram_cell[     668] = 32'h720b12bd;
    ram_cell[     669] = 32'ha7d7465d;
    ram_cell[     670] = 32'hc73ad6ce;
    ram_cell[     671] = 32'h423e5ca6;
    ram_cell[     672] = 32'h47c86971;
    ram_cell[     673] = 32'h14dfc244;
    ram_cell[     674] = 32'h17bdc516;
    ram_cell[     675] = 32'h937e84ce;
    ram_cell[     676] = 32'hb036154b;
    ram_cell[     677] = 32'h1af438f2;
    ram_cell[     678] = 32'h632c90ea;
    ram_cell[     679] = 32'h38100ad8;
    ram_cell[     680] = 32'he829f068;
    ram_cell[     681] = 32'hff569e48;
    ram_cell[     682] = 32'hccae7f93;
    ram_cell[     683] = 32'hab23eebc;
    ram_cell[     684] = 32'heb570410;
    ram_cell[     685] = 32'h34cfe9ec;
    ram_cell[     686] = 32'he35d4905;
    ram_cell[     687] = 32'haa054e45;
    ram_cell[     688] = 32'hbed926b1;
    ram_cell[     689] = 32'h81d8ffd8;
    ram_cell[     690] = 32'hd87bef35;
    ram_cell[     691] = 32'hd707a72f;
    ram_cell[     692] = 32'h014d2a06;
    ram_cell[     693] = 32'hdaee13d2;
    ram_cell[     694] = 32'hc1262747;
    ram_cell[     695] = 32'haf6c4513;
    ram_cell[     696] = 32'h3b60af01;
    ram_cell[     697] = 32'hc9aa2d46;
    ram_cell[     698] = 32'h92c236bd;
    ram_cell[     699] = 32'hc3244b3d;
    ram_cell[     700] = 32'hb974b27a;
    ram_cell[     701] = 32'h4cd2928e;
    ram_cell[     702] = 32'ha73ab0df;
    ram_cell[     703] = 32'hb2f9bf99;
    ram_cell[     704] = 32'he154ed09;
    ram_cell[     705] = 32'hccd52890;
    ram_cell[     706] = 32'had07e58a;
    ram_cell[     707] = 32'h4e92df74;
    ram_cell[     708] = 32'h70ebff0c;
    ram_cell[     709] = 32'h4f6a4c7e;
    ram_cell[     710] = 32'h808f5529;
    ram_cell[     711] = 32'h52b04034;
    ram_cell[     712] = 32'h99a9d992;
    ram_cell[     713] = 32'h95b2774e;
    ram_cell[     714] = 32'h488b6835;
    ram_cell[     715] = 32'h2bd27d05;
    ram_cell[     716] = 32'he71f04cb;
    ram_cell[     717] = 32'hcba2924b;
    ram_cell[     718] = 32'hfe1c9b6d;
    ram_cell[     719] = 32'ha364acea;
    ram_cell[     720] = 32'hd3cbd12e;
    ram_cell[     721] = 32'hf7b01691;
    ram_cell[     722] = 32'hbdfdab57;
    ram_cell[     723] = 32'hf25f97e4;
    ram_cell[     724] = 32'h07b163b8;
    ram_cell[     725] = 32'h1fd69c70;
    ram_cell[     726] = 32'hc6392b33;
    ram_cell[     727] = 32'hd4d78dc5;
    ram_cell[     728] = 32'he374eb01;
    ram_cell[     729] = 32'h6e5e04ce;
    ram_cell[     730] = 32'h503b4f89;
    ram_cell[     731] = 32'h2d0a9806;
    ram_cell[     732] = 32'ha0c0bdca;
    ram_cell[     733] = 32'h1a323a39;
    ram_cell[     734] = 32'h9e1e181a;
    ram_cell[     735] = 32'h14c11a84;
    ram_cell[     736] = 32'h3b2f0460;
    ram_cell[     737] = 32'h920c062a;
    ram_cell[     738] = 32'ha1bb0ff8;
    ram_cell[     739] = 32'h1949bdfb;
    ram_cell[     740] = 32'h6cff5b85;
    ram_cell[     741] = 32'h37a8c557;
    ram_cell[     742] = 32'he86892c9;
    ram_cell[     743] = 32'h029dd2f2;
    ram_cell[     744] = 32'h74eb079a;
    ram_cell[     745] = 32'hda91f500;
    ram_cell[     746] = 32'ha6959fa7;
    ram_cell[     747] = 32'h64182926;
    ram_cell[     748] = 32'h791c4510;
    ram_cell[     749] = 32'h341ee2d4;
    ram_cell[     750] = 32'heba202a4;
    ram_cell[     751] = 32'h1542b73c;
    ram_cell[     752] = 32'h3a22b217;
    ram_cell[     753] = 32'h7af6bb14;
    ram_cell[     754] = 32'h880df99e;
    ram_cell[     755] = 32'h1c75ce7b;
    ram_cell[     756] = 32'h4685e851;
    ram_cell[     757] = 32'h252089bc;
    ram_cell[     758] = 32'hf0d22981;
    ram_cell[     759] = 32'hd1f7c97c;
    ram_cell[     760] = 32'hf465e30b;
    ram_cell[     761] = 32'h3d32fb43;
    ram_cell[     762] = 32'h67cefbb7;
    ram_cell[     763] = 32'h8abf65e6;
    ram_cell[     764] = 32'he2e30a84;
    ram_cell[     765] = 32'h3c0f1e1c;
    ram_cell[     766] = 32'hf6073fe7;
    ram_cell[     767] = 32'hce807031;
end

endmodule

