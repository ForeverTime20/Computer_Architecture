
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h22c0fb88;
    ram_cell[       1] = 32'h0;  // 32'h5c27a0fe;
    ram_cell[       2] = 32'h0;  // 32'hfdf8e687;
    ram_cell[       3] = 32'h0;  // 32'h5d1faa5e;
    ram_cell[       4] = 32'h0;  // 32'h61f8c361;
    ram_cell[       5] = 32'h0;  // 32'h73e13f39;
    ram_cell[       6] = 32'h0;  // 32'h7d463dbd;
    ram_cell[       7] = 32'h0;  // 32'h876086e4;
    ram_cell[       8] = 32'h0;  // 32'hcbbca4fa;
    ram_cell[       9] = 32'h0;  // 32'h1fb65190;
    ram_cell[      10] = 32'h0;  // 32'h4a7d6f50;
    ram_cell[      11] = 32'h0;  // 32'hbb2eab67;
    ram_cell[      12] = 32'h0;  // 32'hc1c82d72;
    ram_cell[      13] = 32'h0;  // 32'hd3c54e8a;
    ram_cell[      14] = 32'h0;  // 32'h692a75dc;
    ram_cell[      15] = 32'h0;  // 32'h7f29d9f6;
    ram_cell[      16] = 32'h0;  // 32'h05e7d986;
    ram_cell[      17] = 32'h0;  // 32'hf65cb142;
    ram_cell[      18] = 32'h0;  // 32'hefa13237;
    ram_cell[      19] = 32'h0;  // 32'he7523b54;
    ram_cell[      20] = 32'h0;  // 32'h34f434b6;
    ram_cell[      21] = 32'h0;  // 32'h16e751fe;
    ram_cell[      22] = 32'h0;  // 32'hf4336beb;
    ram_cell[      23] = 32'h0;  // 32'h62809772;
    ram_cell[      24] = 32'h0;  // 32'hb1a50856;
    ram_cell[      25] = 32'h0;  // 32'h3d259baa;
    ram_cell[      26] = 32'h0;  // 32'hb5eb2d21;
    ram_cell[      27] = 32'h0;  // 32'h81bf39c2;
    ram_cell[      28] = 32'h0;  // 32'hebe6357b;
    ram_cell[      29] = 32'h0;  // 32'h39bc17c2;
    ram_cell[      30] = 32'h0;  // 32'hd22cf928;
    ram_cell[      31] = 32'h0;  // 32'h9d4bdd3b;
    ram_cell[      32] = 32'h0;  // 32'h3d682f40;
    ram_cell[      33] = 32'h0;  // 32'hda110cf5;
    ram_cell[      34] = 32'h0;  // 32'h3101e538;
    ram_cell[      35] = 32'h0;  // 32'hfe99dc63;
    ram_cell[      36] = 32'h0;  // 32'ha372062a;
    ram_cell[      37] = 32'h0;  // 32'hb21322b8;
    ram_cell[      38] = 32'h0;  // 32'h2e20a8c7;
    ram_cell[      39] = 32'h0;  // 32'h2a41144a;
    ram_cell[      40] = 32'h0;  // 32'hed4c0157;
    ram_cell[      41] = 32'h0;  // 32'h78d1c015;
    ram_cell[      42] = 32'h0;  // 32'hf82e44a4;
    ram_cell[      43] = 32'h0;  // 32'h04bc2d7f;
    ram_cell[      44] = 32'h0;  // 32'h00e840ec;
    ram_cell[      45] = 32'h0;  // 32'h092b884b;
    ram_cell[      46] = 32'h0;  // 32'he2915eaa;
    ram_cell[      47] = 32'h0;  // 32'h1eae80e9;
    ram_cell[      48] = 32'h0;  // 32'h34504868;
    ram_cell[      49] = 32'h0;  // 32'h0551a683;
    ram_cell[      50] = 32'h0;  // 32'h9ed82827;
    ram_cell[      51] = 32'h0;  // 32'hdda1ac2c;
    ram_cell[      52] = 32'h0;  // 32'h32e7ba11;
    ram_cell[      53] = 32'h0;  // 32'hbcf81884;
    ram_cell[      54] = 32'h0;  // 32'h655bc98a;
    ram_cell[      55] = 32'h0;  // 32'h65a3669f;
    ram_cell[      56] = 32'h0;  // 32'h0240be1c;
    ram_cell[      57] = 32'h0;  // 32'h081e5173;
    ram_cell[      58] = 32'h0;  // 32'he2eb6532;
    ram_cell[      59] = 32'h0;  // 32'hd0f5614e;
    ram_cell[      60] = 32'h0;  // 32'h68c62d58;
    ram_cell[      61] = 32'h0;  // 32'h967e7150;
    ram_cell[      62] = 32'h0;  // 32'h3dac5da3;
    ram_cell[      63] = 32'h0;  // 32'h85b9d21b;
    ram_cell[      64] = 32'h0;  // 32'h8d51aad5;
    ram_cell[      65] = 32'h0;  // 32'h67fd0763;
    ram_cell[      66] = 32'h0;  // 32'hf38e24b9;
    ram_cell[      67] = 32'h0;  // 32'h6997aac3;
    ram_cell[      68] = 32'h0;  // 32'h764b77d5;
    ram_cell[      69] = 32'h0;  // 32'hfb7e7604;
    ram_cell[      70] = 32'h0;  // 32'h8ae3e9d3;
    ram_cell[      71] = 32'h0;  // 32'h7f72d3bb;
    ram_cell[      72] = 32'h0;  // 32'h26bae93c;
    ram_cell[      73] = 32'h0;  // 32'h73e85251;
    ram_cell[      74] = 32'h0;  // 32'hd2283126;
    ram_cell[      75] = 32'h0;  // 32'ha8be4f98;
    ram_cell[      76] = 32'h0;  // 32'h4c35b0bb;
    ram_cell[      77] = 32'h0;  // 32'hb68fd04c;
    ram_cell[      78] = 32'h0;  // 32'hff7018e7;
    ram_cell[      79] = 32'h0;  // 32'h5a590640;
    ram_cell[      80] = 32'h0;  // 32'h1fd0443a;
    ram_cell[      81] = 32'h0;  // 32'h142a2b87;
    ram_cell[      82] = 32'h0;  // 32'h7bf04d99;
    ram_cell[      83] = 32'h0;  // 32'h52e7a2c1;
    ram_cell[      84] = 32'h0;  // 32'h428eb732;
    ram_cell[      85] = 32'h0;  // 32'h17efe461;
    ram_cell[      86] = 32'h0;  // 32'h29e46c5f;
    ram_cell[      87] = 32'h0;  // 32'h3c36a226;
    ram_cell[      88] = 32'h0;  // 32'h51ce0dfd;
    ram_cell[      89] = 32'h0;  // 32'h44f7d43e;
    ram_cell[      90] = 32'h0;  // 32'h211bda7d;
    ram_cell[      91] = 32'h0;  // 32'h3b29f035;
    ram_cell[      92] = 32'h0;  // 32'h89da767e;
    ram_cell[      93] = 32'h0;  // 32'hea9ecd8b;
    ram_cell[      94] = 32'h0;  // 32'h65942ccd;
    ram_cell[      95] = 32'h0;  // 32'hd7911ca3;
    ram_cell[      96] = 32'h0;  // 32'h1c2ab6b9;
    ram_cell[      97] = 32'h0;  // 32'h530aa32e;
    ram_cell[      98] = 32'h0;  // 32'hc6b2a996;
    ram_cell[      99] = 32'h0;  // 32'h115e1e08;
    ram_cell[     100] = 32'h0;  // 32'h06460c95;
    ram_cell[     101] = 32'h0;  // 32'hcf783c21;
    ram_cell[     102] = 32'h0;  // 32'h225aff4f;
    ram_cell[     103] = 32'h0;  // 32'h5135ffcb;
    ram_cell[     104] = 32'h0;  // 32'he877de2b;
    ram_cell[     105] = 32'h0;  // 32'hd1bdc27b;
    ram_cell[     106] = 32'h0;  // 32'hfaa1679d;
    ram_cell[     107] = 32'h0;  // 32'he6617b8b;
    ram_cell[     108] = 32'h0;  // 32'hdb8bf9ee;
    ram_cell[     109] = 32'h0;  // 32'h2c4cda33;
    ram_cell[     110] = 32'h0;  // 32'h8f30d794;
    ram_cell[     111] = 32'h0;  // 32'hce3ad14d;
    ram_cell[     112] = 32'h0;  // 32'hf8106d3d;
    ram_cell[     113] = 32'h0;  // 32'he3a4bb46;
    ram_cell[     114] = 32'h0;  // 32'h7342df97;
    ram_cell[     115] = 32'h0;  // 32'hb25eff38;
    ram_cell[     116] = 32'h0;  // 32'h1a58090e;
    ram_cell[     117] = 32'h0;  // 32'hc75a4bf1;
    ram_cell[     118] = 32'h0;  // 32'h902cdca0;
    ram_cell[     119] = 32'h0;  // 32'h7240f822;
    ram_cell[     120] = 32'h0;  // 32'h4d1974ec;
    ram_cell[     121] = 32'h0;  // 32'h4f11244b;
    ram_cell[     122] = 32'h0;  // 32'hfe60af93;
    ram_cell[     123] = 32'h0;  // 32'h60c82dce;
    ram_cell[     124] = 32'h0;  // 32'h8eb3fb82;
    ram_cell[     125] = 32'h0;  // 32'h96da51ce;
    ram_cell[     126] = 32'h0;  // 32'h45972f42;
    ram_cell[     127] = 32'h0;  // 32'hcd0d7ca4;
    ram_cell[     128] = 32'h0;  // 32'h7d725cfa;
    ram_cell[     129] = 32'h0;  // 32'h5db3fc13;
    ram_cell[     130] = 32'h0;  // 32'h536c5fe9;
    ram_cell[     131] = 32'h0;  // 32'h48ac1a9e;
    ram_cell[     132] = 32'h0;  // 32'h3e5c4e1f;
    ram_cell[     133] = 32'h0;  // 32'hc7de412b;
    ram_cell[     134] = 32'h0;  // 32'hdb01ca62;
    ram_cell[     135] = 32'h0;  // 32'h93257fde;
    ram_cell[     136] = 32'h0;  // 32'h486ce9b6;
    ram_cell[     137] = 32'h0;  // 32'hdce0ee5f;
    ram_cell[     138] = 32'h0;  // 32'hc5bbccb7;
    ram_cell[     139] = 32'h0;  // 32'hc8aab303;
    ram_cell[     140] = 32'h0;  // 32'h1e09f6e8;
    ram_cell[     141] = 32'h0;  // 32'h522ae21e;
    ram_cell[     142] = 32'h0;  // 32'ha67efb00;
    ram_cell[     143] = 32'h0;  // 32'hb1b8c92d;
    ram_cell[     144] = 32'h0;  // 32'he264513b;
    ram_cell[     145] = 32'h0;  // 32'h333e8e95;
    ram_cell[     146] = 32'h0;  // 32'h4b5e5392;
    ram_cell[     147] = 32'h0;  // 32'h9e5ee7a9;
    ram_cell[     148] = 32'h0;  // 32'h94d92561;
    ram_cell[     149] = 32'h0;  // 32'he2140e22;
    ram_cell[     150] = 32'h0;  // 32'hb0ace7b7;
    ram_cell[     151] = 32'h0;  // 32'hef141d9b;
    ram_cell[     152] = 32'h0;  // 32'hae523b67;
    ram_cell[     153] = 32'h0;  // 32'h50e79ed4;
    ram_cell[     154] = 32'h0;  // 32'he5d32f28;
    ram_cell[     155] = 32'h0;  // 32'ha2f38854;
    ram_cell[     156] = 32'h0;  // 32'h02532f3f;
    ram_cell[     157] = 32'h0;  // 32'hd482c4d0;
    ram_cell[     158] = 32'h0;  // 32'heea94300;
    ram_cell[     159] = 32'h0;  // 32'h65008a84;
    ram_cell[     160] = 32'h0;  // 32'he36225d1;
    ram_cell[     161] = 32'h0;  // 32'hff165c83;
    ram_cell[     162] = 32'h0;  // 32'h88bf87b5;
    ram_cell[     163] = 32'h0;  // 32'hbdd52a3c;
    ram_cell[     164] = 32'h0;  // 32'hd87c3700;
    ram_cell[     165] = 32'h0;  // 32'h87422e6a;
    ram_cell[     166] = 32'h0;  // 32'h289d1bbc;
    ram_cell[     167] = 32'h0;  // 32'h790eec33;
    ram_cell[     168] = 32'h0;  // 32'h03c8fc5f;
    ram_cell[     169] = 32'h0;  // 32'hb170f24f;
    ram_cell[     170] = 32'h0;  // 32'h436614c3;
    ram_cell[     171] = 32'h0;  // 32'hfc1332d6;
    ram_cell[     172] = 32'h0;  // 32'h0f6126d2;
    ram_cell[     173] = 32'h0;  // 32'h6c45a8cd;
    ram_cell[     174] = 32'h0;  // 32'h4c7620b1;
    ram_cell[     175] = 32'h0;  // 32'hc34e185d;
    ram_cell[     176] = 32'h0;  // 32'h33496c21;
    ram_cell[     177] = 32'h0;  // 32'he4d304ae;
    ram_cell[     178] = 32'h0;  // 32'h3fca51a6;
    ram_cell[     179] = 32'h0;  // 32'h170cced6;
    ram_cell[     180] = 32'h0;  // 32'h75d6102f;
    ram_cell[     181] = 32'h0;  // 32'h7ef030a8;
    ram_cell[     182] = 32'h0;  // 32'h5a45c9d4;
    ram_cell[     183] = 32'h0;  // 32'h32bea0c5;
    ram_cell[     184] = 32'h0;  // 32'ha1c7ad82;
    ram_cell[     185] = 32'h0;  // 32'he4bdcf1c;
    ram_cell[     186] = 32'h0;  // 32'h97a386e4;
    ram_cell[     187] = 32'h0;  // 32'h49a27d09;
    ram_cell[     188] = 32'h0;  // 32'h2d3f2b1f;
    ram_cell[     189] = 32'h0;  // 32'h070c9fbd;
    ram_cell[     190] = 32'h0;  // 32'h553abcf8;
    ram_cell[     191] = 32'h0;  // 32'h07e5e742;
    ram_cell[     192] = 32'h0;  // 32'h438454e0;
    ram_cell[     193] = 32'h0;  // 32'h1cc63398;
    ram_cell[     194] = 32'h0;  // 32'h32976b59;
    ram_cell[     195] = 32'h0;  // 32'h24e628ff;
    ram_cell[     196] = 32'h0;  // 32'h897c7a3c;
    ram_cell[     197] = 32'h0;  // 32'h6011c958;
    ram_cell[     198] = 32'h0;  // 32'h3df0f3e9;
    ram_cell[     199] = 32'h0;  // 32'h356cd4e1;
    ram_cell[     200] = 32'h0;  // 32'hfe3e7d6b;
    ram_cell[     201] = 32'h0;  // 32'h3a3ffc53;
    ram_cell[     202] = 32'h0;  // 32'h1f2a0cd7;
    ram_cell[     203] = 32'h0;  // 32'h77d9a3e3;
    ram_cell[     204] = 32'h0;  // 32'h00d003e6;
    ram_cell[     205] = 32'h0;  // 32'h8e4e29f4;
    ram_cell[     206] = 32'h0;  // 32'h721924dc;
    ram_cell[     207] = 32'h0;  // 32'hb578a7ad;
    ram_cell[     208] = 32'h0;  // 32'h74526d80;
    ram_cell[     209] = 32'h0;  // 32'hbd20ce63;
    ram_cell[     210] = 32'h0;  // 32'hf2f83de6;
    ram_cell[     211] = 32'h0;  // 32'h25169451;
    ram_cell[     212] = 32'h0;  // 32'hbfed80bd;
    ram_cell[     213] = 32'h0;  // 32'hd89248e0;
    ram_cell[     214] = 32'h0;  // 32'h94bb55f3;
    ram_cell[     215] = 32'h0;  // 32'h519f3891;
    ram_cell[     216] = 32'h0;  // 32'h8f11105b;
    ram_cell[     217] = 32'h0;  // 32'haf9e7888;
    ram_cell[     218] = 32'h0;  // 32'hc56b61c2;
    ram_cell[     219] = 32'h0;  // 32'h0dff7d52;
    ram_cell[     220] = 32'h0;  // 32'hb2effc30;
    ram_cell[     221] = 32'h0;  // 32'h0f4e477d;
    ram_cell[     222] = 32'h0;  // 32'h5e7fa4e7;
    ram_cell[     223] = 32'h0;  // 32'h8e27911c;
    ram_cell[     224] = 32'h0;  // 32'h5f58d585;
    ram_cell[     225] = 32'h0;  // 32'hf3692a1c;
    ram_cell[     226] = 32'h0;  // 32'h5abacf02;
    ram_cell[     227] = 32'h0;  // 32'hf710fc90;
    ram_cell[     228] = 32'h0;  // 32'h448e0bee;
    ram_cell[     229] = 32'h0;  // 32'h264321e0;
    ram_cell[     230] = 32'h0;  // 32'h2f8f0a0b;
    ram_cell[     231] = 32'h0;  // 32'ha399825b;
    ram_cell[     232] = 32'h0;  // 32'h42b61113;
    ram_cell[     233] = 32'h0;  // 32'h6a18d6de;
    ram_cell[     234] = 32'h0;  // 32'hcf473c5f;
    ram_cell[     235] = 32'h0;  // 32'hc752176c;
    ram_cell[     236] = 32'h0;  // 32'he1bbbcb9;
    ram_cell[     237] = 32'h0;  // 32'h9cce8a34;
    ram_cell[     238] = 32'h0;  // 32'h003c697c;
    ram_cell[     239] = 32'h0;  // 32'hfa95fec6;
    ram_cell[     240] = 32'h0;  // 32'hea6a78e2;
    ram_cell[     241] = 32'h0;  // 32'h3a7422b8;
    ram_cell[     242] = 32'h0;  // 32'h28f6b3a3;
    ram_cell[     243] = 32'h0;  // 32'h0bb0f1e5;
    ram_cell[     244] = 32'h0;  // 32'ha1aafb5e;
    ram_cell[     245] = 32'h0;  // 32'h8c46b4ba;
    ram_cell[     246] = 32'h0;  // 32'h07c85b1d;
    ram_cell[     247] = 32'h0;  // 32'h50977f8b;
    ram_cell[     248] = 32'h0;  // 32'h249c5133;
    ram_cell[     249] = 32'h0;  // 32'h683e9fd1;
    ram_cell[     250] = 32'h0;  // 32'h8575b96b;
    ram_cell[     251] = 32'h0;  // 32'h4a06dfd1;
    ram_cell[     252] = 32'h0;  // 32'h6f4fcc65;
    ram_cell[     253] = 32'h0;  // 32'he980eead;
    ram_cell[     254] = 32'h0;  // 32'h96ac6da6;
    ram_cell[     255] = 32'h0;  // 32'hc9ec309c;
    // src matrix A
    ram_cell[     256] = 32'h5e96b1d9;
    ram_cell[     257] = 32'hbf79f3fc;
    ram_cell[     258] = 32'he6150ccb;
    ram_cell[     259] = 32'he39282df;
    ram_cell[     260] = 32'hc34b56e8;
    ram_cell[     261] = 32'h24823ba1;
    ram_cell[     262] = 32'h8120a4e0;
    ram_cell[     263] = 32'h8df4751d;
    ram_cell[     264] = 32'hbdbda1d7;
    ram_cell[     265] = 32'h2313b1bc;
    ram_cell[     266] = 32'h5dbce577;
    ram_cell[     267] = 32'hf7b961ef;
    ram_cell[     268] = 32'h2d31d570;
    ram_cell[     269] = 32'hbd2de2cb;
    ram_cell[     270] = 32'ha516177e;
    ram_cell[     271] = 32'h43c02406;
    ram_cell[     272] = 32'hb963f754;
    ram_cell[     273] = 32'h40f32c3d;
    ram_cell[     274] = 32'h30648d1e;
    ram_cell[     275] = 32'h03c9467e;
    ram_cell[     276] = 32'h838648d0;
    ram_cell[     277] = 32'haa3ac2f6;
    ram_cell[     278] = 32'h8f1f90da;
    ram_cell[     279] = 32'haeba4ed8;
    ram_cell[     280] = 32'h2ff7e85d;
    ram_cell[     281] = 32'h6dff73dd;
    ram_cell[     282] = 32'h0b66de28;
    ram_cell[     283] = 32'h7f2c97ac;
    ram_cell[     284] = 32'h4a71b315;
    ram_cell[     285] = 32'h22b9f1cf;
    ram_cell[     286] = 32'h5864462c;
    ram_cell[     287] = 32'h8124891c;
    ram_cell[     288] = 32'hb091eb9e;
    ram_cell[     289] = 32'h2817bc1d;
    ram_cell[     290] = 32'h488817fd;
    ram_cell[     291] = 32'hfeae7f53;
    ram_cell[     292] = 32'h9770315b;
    ram_cell[     293] = 32'h12bbcd0f;
    ram_cell[     294] = 32'hf2d4555c;
    ram_cell[     295] = 32'h3a4a486c;
    ram_cell[     296] = 32'hed5773cf;
    ram_cell[     297] = 32'h8e6e493e;
    ram_cell[     298] = 32'hd776f1fd;
    ram_cell[     299] = 32'h5f7d0af5;
    ram_cell[     300] = 32'h3711ed5f;
    ram_cell[     301] = 32'ha5b08d08;
    ram_cell[     302] = 32'hffe58c99;
    ram_cell[     303] = 32'h449e40ff;
    ram_cell[     304] = 32'h45e5fb17;
    ram_cell[     305] = 32'h1f7ff452;
    ram_cell[     306] = 32'h08173ddd;
    ram_cell[     307] = 32'haa761eeb;
    ram_cell[     308] = 32'he53e7811;
    ram_cell[     309] = 32'h4f97879c;
    ram_cell[     310] = 32'h0a25d7dc;
    ram_cell[     311] = 32'ha8c308a1;
    ram_cell[     312] = 32'hd7645efb;
    ram_cell[     313] = 32'hc1892c74;
    ram_cell[     314] = 32'he89270a9;
    ram_cell[     315] = 32'h65321929;
    ram_cell[     316] = 32'hcf81545f;
    ram_cell[     317] = 32'hb2cd48a1;
    ram_cell[     318] = 32'h6c62446b;
    ram_cell[     319] = 32'h002a82d8;
    ram_cell[     320] = 32'heabe80ba;
    ram_cell[     321] = 32'h7617ea05;
    ram_cell[     322] = 32'h3e4418df;
    ram_cell[     323] = 32'h99bc979c;
    ram_cell[     324] = 32'hbe1465aa;
    ram_cell[     325] = 32'h35dbe397;
    ram_cell[     326] = 32'hc37e1526;
    ram_cell[     327] = 32'h3c637d57;
    ram_cell[     328] = 32'h8d4c9d1e;
    ram_cell[     329] = 32'h05d803df;
    ram_cell[     330] = 32'h05bece26;
    ram_cell[     331] = 32'h8d8fb728;
    ram_cell[     332] = 32'hd0f4e7e8;
    ram_cell[     333] = 32'h933da6ed;
    ram_cell[     334] = 32'h766f322b;
    ram_cell[     335] = 32'hb74a7225;
    ram_cell[     336] = 32'h79afa417;
    ram_cell[     337] = 32'h4060fedf;
    ram_cell[     338] = 32'h3ea45278;
    ram_cell[     339] = 32'hb279a8da;
    ram_cell[     340] = 32'hdc6961fe;
    ram_cell[     341] = 32'h3cadc2dc;
    ram_cell[     342] = 32'h9119f551;
    ram_cell[     343] = 32'h717b595c;
    ram_cell[     344] = 32'h0a1d7158;
    ram_cell[     345] = 32'h55faabf0;
    ram_cell[     346] = 32'h9adfd8ee;
    ram_cell[     347] = 32'h7064a9fe;
    ram_cell[     348] = 32'he75b07e8;
    ram_cell[     349] = 32'h200042de;
    ram_cell[     350] = 32'hebfba297;
    ram_cell[     351] = 32'he9c948db;
    ram_cell[     352] = 32'hb58bcaa6;
    ram_cell[     353] = 32'hb8c0cbe9;
    ram_cell[     354] = 32'hf4073756;
    ram_cell[     355] = 32'h38a20fab;
    ram_cell[     356] = 32'h15b65e7e;
    ram_cell[     357] = 32'h041dd36d;
    ram_cell[     358] = 32'h36a9abb1;
    ram_cell[     359] = 32'h17818695;
    ram_cell[     360] = 32'h6ec3741e;
    ram_cell[     361] = 32'h75ad2bda;
    ram_cell[     362] = 32'hd3666f14;
    ram_cell[     363] = 32'hec5f980a;
    ram_cell[     364] = 32'h7cfb3ea8;
    ram_cell[     365] = 32'h9f0943c2;
    ram_cell[     366] = 32'hca0fec99;
    ram_cell[     367] = 32'h2959023e;
    ram_cell[     368] = 32'h4c8371de;
    ram_cell[     369] = 32'h56aed332;
    ram_cell[     370] = 32'he6e4794d;
    ram_cell[     371] = 32'h3fda8b46;
    ram_cell[     372] = 32'h814a179a;
    ram_cell[     373] = 32'h24105729;
    ram_cell[     374] = 32'hcab345b7;
    ram_cell[     375] = 32'hccbe0216;
    ram_cell[     376] = 32'he78ae45f;
    ram_cell[     377] = 32'ha642ed37;
    ram_cell[     378] = 32'h444f0718;
    ram_cell[     379] = 32'h3ffc21b7;
    ram_cell[     380] = 32'haf68d40e;
    ram_cell[     381] = 32'h600c0337;
    ram_cell[     382] = 32'hc2bd1217;
    ram_cell[     383] = 32'h57c19a39;
    ram_cell[     384] = 32'h51bea14c;
    ram_cell[     385] = 32'h6e70149e;
    ram_cell[     386] = 32'h0d2fb750;
    ram_cell[     387] = 32'ha6701a8d;
    ram_cell[     388] = 32'h368bfc6e;
    ram_cell[     389] = 32'h2e923d28;
    ram_cell[     390] = 32'haa6be133;
    ram_cell[     391] = 32'h6608c108;
    ram_cell[     392] = 32'he5922ada;
    ram_cell[     393] = 32'h97928eb9;
    ram_cell[     394] = 32'h81c4c204;
    ram_cell[     395] = 32'h84b2e0ac;
    ram_cell[     396] = 32'h5776d355;
    ram_cell[     397] = 32'h4ee30066;
    ram_cell[     398] = 32'h9f211bf8;
    ram_cell[     399] = 32'h868a534c;
    ram_cell[     400] = 32'hef53badb;
    ram_cell[     401] = 32'h474890df;
    ram_cell[     402] = 32'h155fe414;
    ram_cell[     403] = 32'h1c579827;
    ram_cell[     404] = 32'h499529d4;
    ram_cell[     405] = 32'h1c7e3e82;
    ram_cell[     406] = 32'h258c247f;
    ram_cell[     407] = 32'he1bb62aa;
    ram_cell[     408] = 32'hc771ef50;
    ram_cell[     409] = 32'h79c49fd7;
    ram_cell[     410] = 32'h5de75967;
    ram_cell[     411] = 32'hc1a488e0;
    ram_cell[     412] = 32'h7bd20e85;
    ram_cell[     413] = 32'hc97671e7;
    ram_cell[     414] = 32'he3ce9561;
    ram_cell[     415] = 32'h4be43da5;
    ram_cell[     416] = 32'h0ef35784;
    ram_cell[     417] = 32'h16031f53;
    ram_cell[     418] = 32'h2db9ef14;
    ram_cell[     419] = 32'h9d7dbee7;
    ram_cell[     420] = 32'h7bacbc37;
    ram_cell[     421] = 32'hc6eb8807;
    ram_cell[     422] = 32'h2e53478d;
    ram_cell[     423] = 32'h985c3f2b;
    ram_cell[     424] = 32'hda1b21c4;
    ram_cell[     425] = 32'h2f636b68;
    ram_cell[     426] = 32'h8c70bfd5;
    ram_cell[     427] = 32'h193c0b58;
    ram_cell[     428] = 32'h7d8a9105;
    ram_cell[     429] = 32'h7e4a2594;
    ram_cell[     430] = 32'hfd8e0df5;
    ram_cell[     431] = 32'hc07693bc;
    ram_cell[     432] = 32'h6369b89d;
    ram_cell[     433] = 32'h53829cee;
    ram_cell[     434] = 32'hfacc0f92;
    ram_cell[     435] = 32'h6e03bba9;
    ram_cell[     436] = 32'h62448036;
    ram_cell[     437] = 32'h2ae98918;
    ram_cell[     438] = 32'h3f5760bb;
    ram_cell[     439] = 32'h58b32e2b;
    ram_cell[     440] = 32'h0637ea4f;
    ram_cell[     441] = 32'hb1a2d6c0;
    ram_cell[     442] = 32'h8a61b089;
    ram_cell[     443] = 32'h862eee10;
    ram_cell[     444] = 32'h3246057b;
    ram_cell[     445] = 32'h31fd6f08;
    ram_cell[     446] = 32'h85fae2f8;
    ram_cell[     447] = 32'hab64f759;
    ram_cell[     448] = 32'h8103a411;
    ram_cell[     449] = 32'h70573eed;
    ram_cell[     450] = 32'h63007acd;
    ram_cell[     451] = 32'h2b6316c9;
    ram_cell[     452] = 32'hcde5b4b3;
    ram_cell[     453] = 32'he24763fd;
    ram_cell[     454] = 32'h038172b0;
    ram_cell[     455] = 32'h2e184087;
    ram_cell[     456] = 32'h2692fd30;
    ram_cell[     457] = 32'h345d3825;
    ram_cell[     458] = 32'hb1aefdd7;
    ram_cell[     459] = 32'h9b532574;
    ram_cell[     460] = 32'ha2b72d6c;
    ram_cell[     461] = 32'h28fe7ddc;
    ram_cell[     462] = 32'h8890c813;
    ram_cell[     463] = 32'he753835f;
    ram_cell[     464] = 32'hcceb6c11;
    ram_cell[     465] = 32'h885d0b83;
    ram_cell[     466] = 32'ha2b98e60;
    ram_cell[     467] = 32'h41716922;
    ram_cell[     468] = 32'h39d9e117;
    ram_cell[     469] = 32'hec778e9c;
    ram_cell[     470] = 32'h6e4f9aa3;
    ram_cell[     471] = 32'h9c698f7c;
    ram_cell[     472] = 32'h8caeb067;
    ram_cell[     473] = 32'hf1d9c9e5;
    ram_cell[     474] = 32'h09b7efc5;
    ram_cell[     475] = 32'h48a08aa1;
    ram_cell[     476] = 32'h564d40b6;
    ram_cell[     477] = 32'h0a4c4963;
    ram_cell[     478] = 32'h8c20209c;
    ram_cell[     479] = 32'h215aba69;
    ram_cell[     480] = 32'h1cf15b95;
    ram_cell[     481] = 32'h3e39f654;
    ram_cell[     482] = 32'h333fb713;
    ram_cell[     483] = 32'he3cc5df0;
    ram_cell[     484] = 32'h6a6f7e3c;
    ram_cell[     485] = 32'he2615e6c;
    ram_cell[     486] = 32'hf75f309f;
    ram_cell[     487] = 32'h493aa054;
    ram_cell[     488] = 32'h91751759;
    ram_cell[     489] = 32'h90711835;
    ram_cell[     490] = 32'h6fc1329a;
    ram_cell[     491] = 32'ha2f03490;
    ram_cell[     492] = 32'haefb2e35;
    ram_cell[     493] = 32'hbbcb3497;
    ram_cell[     494] = 32'h1d88ffc5;
    ram_cell[     495] = 32'hda2e208f;
    ram_cell[     496] = 32'h328eba57;
    ram_cell[     497] = 32'h8813edb2;
    ram_cell[     498] = 32'h88a52a23;
    ram_cell[     499] = 32'h42b9f210;
    ram_cell[     500] = 32'hb15cf008;
    ram_cell[     501] = 32'hb32e9869;
    ram_cell[     502] = 32'h388fe19d;
    ram_cell[     503] = 32'h3b4df74d;
    ram_cell[     504] = 32'h800f17f7;
    ram_cell[     505] = 32'h41c4e56e;
    ram_cell[     506] = 32'h892599cd;
    ram_cell[     507] = 32'he0cf823b;
    ram_cell[     508] = 32'h2d6fe41b;
    ram_cell[     509] = 32'h74a11e84;
    ram_cell[     510] = 32'hd8b38357;
    ram_cell[     511] = 32'h0e34a14b;
    // src matrix B
    ram_cell[     512] = 32'hf57420ea;
    ram_cell[     513] = 32'h4b848921;
    ram_cell[     514] = 32'h8826f3b9;
    ram_cell[     515] = 32'h4a41a306;
    ram_cell[     516] = 32'h278887db;
    ram_cell[     517] = 32'h37bd7a9a;
    ram_cell[     518] = 32'h320fed8b;
    ram_cell[     519] = 32'h628554df;
    ram_cell[     520] = 32'hc4b15bc5;
    ram_cell[     521] = 32'hfb852222;
    ram_cell[     522] = 32'hea45b16e;
    ram_cell[     523] = 32'h1de7d0c1;
    ram_cell[     524] = 32'h873b9c47;
    ram_cell[     525] = 32'h1a9bf0dd;
    ram_cell[     526] = 32'h9e6fa4a3;
    ram_cell[     527] = 32'hc4dfdabc;
    ram_cell[     528] = 32'he733b8df;
    ram_cell[     529] = 32'hdacfec29;
    ram_cell[     530] = 32'hded1fff2;
    ram_cell[     531] = 32'hb1533312;
    ram_cell[     532] = 32'he6cb395f;
    ram_cell[     533] = 32'h3e7c90c9;
    ram_cell[     534] = 32'hefc70e6c;
    ram_cell[     535] = 32'h2c2491df;
    ram_cell[     536] = 32'hc9dc6d1d;
    ram_cell[     537] = 32'h8d93643f;
    ram_cell[     538] = 32'h7a168191;
    ram_cell[     539] = 32'h85f979f9;
    ram_cell[     540] = 32'h11b53684;
    ram_cell[     541] = 32'he6461e26;
    ram_cell[     542] = 32'h1a1d9dc7;
    ram_cell[     543] = 32'he4a500de;
    ram_cell[     544] = 32'hbab89149;
    ram_cell[     545] = 32'h18d227e5;
    ram_cell[     546] = 32'hc0c541d6;
    ram_cell[     547] = 32'hac1663ad;
    ram_cell[     548] = 32'hc477e88a;
    ram_cell[     549] = 32'hb041f971;
    ram_cell[     550] = 32'h2fdd027b;
    ram_cell[     551] = 32'h588eaa07;
    ram_cell[     552] = 32'h24e7457a;
    ram_cell[     553] = 32'hb70bcde2;
    ram_cell[     554] = 32'he069d549;
    ram_cell[     555] = 32'h99b01f39;
    ram_cell[     556] = 32'h1b72d03a;
    ram_cell[     557] = 32'h9d32ebff;
    ram_cell[     558] = 32'h99bcadc5;
    ram_cell[     559] = 32'h6cda16e8;
    ram_cell[     560] = 32'h69563b5f;
    ram_cell[     561] = 32'h0e6a9575;
    ram_cell[     562] = 32'h1f350143;
    ram_cell[     563] = 32'h4d5ba85f;
    ram_cell[     564] = 32'hae004dfe;
    ram_cell[     565] = 32'hdc4c70e1;
    ram_cell[     566] = 32'h0d47d472;
    ram_cell[     567] = 32'h7ab52cb4;
    ram_cell[     568] = 32'h4f2ac5e4;
    ram_cell[     569] = 32'h2532472c;
    ram_cell[     570] = 32'hb0977cea;
    ram_cell[     571] = 32'hc60a6229;
    ram_cell[     572] = 32'hc8d93ce6;
    ram_cell[     573] = 32'hdfa78d14;
    ram_cell[     574] = 32'h8ae3121d;
    ram_cell[     575] = 32'hb64bdadf;
    ram_cell[     576] = 32'h1383d67f;
    ram_cell[     577] = 32'h5a689470;
    ram_cell[     578] = 32'hef571945;
    ram_cell[     579] = 32'h596fbfdc;
    ram_cell[     580] = 32'hc7258866;
    ram_cell[     581] = 32'h4bd5b84f;
    ram_cell[     582] = 32'h0d8d8d53;
    ram_cell[     583] = 32'h022cd7a7;
    ram_cell[     584] = 32'h6ba34f6b;
    ram_cell[     585] = 32'h027e0ab9;
    ram_cell[     586] = 32'hf1db7df1;
    ram_cell[     587] = 32'h11701449;
    ram_cell[     588] = 32'h2ed0fc3d;
    ram_cell[     589] = 32'h900e018f;
    ram_cell[     590] = 32'h3c0b9c8c;
    ram_cell[     591] = 32'h18c144db;
    ram_cell[     592] = 32'h94deb878;
    ram_cell[     593] = 32'h5c66ad34;
    ram_cell[     594] = 32'h50c982fb;
    ram_cell[     595] = 32'h5bcad16d;
    ram_cell[     596] = 32'h7251f5c0;
    ram_cell[     597] = 32'hee474be3;
    ram_cell[     598] = 32'h54cfcf50;
    ram_cell[     599] = 32'hb3b28d83;
    ram_cell[     600] = 32'hd94d441c;
    ram_cell[     601] = 32'h06b5710e;
    ram_cell[     602] = 32'h25ebb023;
    ram_cell[     603] = 32'h30dbe509;
    ram_cell[     604] = 32'h49474b2b;
    ram_cell[     605] = 32'h8f3c332d;
    ram_cell[     606] = 32'h7e717c92;
    ram_cell[     607] = 32'h4a304ff9;
    ram_cell[     608] = 32'h536394a6;
    ram_cell[     609] = 32'hd1f1b656;
    ram_cell[     610] = 32'h81e14e6b;
    ram_cell[     611] = 32'h5f024785;
    ram_cell[     612] = 32'h13cd8fa0;
    ram_cell[     613] = 32'hd4611b5e;
    ram_cell[     614] = 32'h5edb5e8c;
    ram_cell[     615] = 32'h205ac8ab;
    ram_cell[     616] = 32'h1b65b72f;
    ram_cell[     617] = 32'hd82d12fa;
    ram_cell[     618] = 32'h9e414a9c;
    ram_cell[     619] = 32'h8b3782d0;
    ram_cell[     620] = 32'h1cc4c9f2;
    ram_cell[     621] = 32'hd6cfe35b;
    ram_cell[     622] = 32'he4eb6452;
    ram_cell[     623] = 32'h64903ad5;
    ram_cell[     624] = 32'hee7b8d33;
    ram_cell[     625] = 32'h3906ad84;
    ram_cell[     626] = 32'hbc64aa37;
    ram_cell[     627] = 32'h5b50aff0;
    ram_cell[     628] = 32'h6ccbc38c;
    ram_cell[     629] = 32'h8ce6367d;
    ram_cell[     630] = 32'h468d50f4;
    ram_cell[     631] = 32'h22471933;
    ram_cell[     632] = 32'h77c49308;
    ram_cell[     633] = 32'h9c21fbfc;
    ram_cell[     634] = 32'hccbe33bb;
    ram_cell[     635] = 32'hcd278398;
    ram_cell[     636] = 32'h040c1d1b;
    ram_cell[     637] = 32'hbc19f161;
    ram_cell[     638] = 32'h706a6eb5;
    ram_cell[     639] = 32'hda1b51fa;
    ram_cell[     640] = 32'hfd96b02d;
    ram_cell[     641] = 32'h69572fee;
    ram_cell[     642] = 32'h4eb8d3ab;
    ram_cell[     643] = 32'hd9be3737;
    ram_cell[     644] = 32'h30556a3d;
    ram_cell[     645] = 32'h32fe110b;
    ram_cell[     646] = 32'hd626d52e;
    ram_cell[     647] = 32'hbb2e5293;
    ram_cell[     648] = 32'he1c1db48;
    ram_cell[     649] = 32'h5a77a8f8;
    ram_cell[     650] = 32'h7363110c;
    ram_cell[     651] = 32'h2b36c4aa;
    ram_cell[     652] = 32'he67a7959;
    ram_cell[     653] = 32'h0ad5dcaa;
    ram_cell[     654] = 32'hafe98768;
    ram_cell[     655] = 32'h5a99a629;
    ram_cell[     656] = 32'h7660c468;
    ram_cell[     657] = 32'hbb5bbad5;
    ram_cell[     658] = 32'hc230e9bf;
    ram_cell[     659] = 32'h6e7c4e9c;
    ram_cell[     660] = 32'h31496a93;
    ram_cell[     661] = 32'hd586f4b2;
    ram_cell[     662] = 32'haf732865;
    ram_cell[     663] = 32'h8f12f993;
    ram_cell[     664] = 32'hbe9efc5d;
    ram_cell[     665] = 32'h059670e9;
    ram_cell[     666] = 32'h2683e86f;
    ram_cell[     667] = 32'hbb1e14c7;
    ram_cell[     668] = 32'hd49bcc72;
    ram_cell[     669] = 32'h31977811;
    ram_cell[     670] = 32'h296f5f43;
    ram_cell[     671] = 32'h23fdf218;
    ram_cell[     672] = 32'h2e83a952;
    ram_cell[     673] = 32'h9b08a588;
    ram_cell[     674] = 32'h85a975dc;
    ram_cell[     675] = 32'h33306836;
    ram_cell[     676] = 32'h932235af;
    ram_cell[     677] = 32'h256915c6;
    ram_cell[     678] = 32'h81b1873d;
    ram_cell[     679] = 32'h14929bb9;
    ram_cell[     680] = 32'hb9392acf;
    ram_cell[     681] = 32'h98d197d3;
    ram_cell[     682] = 32'h6a2e7a79;
    ram_cell[     683] = 32'hf555fd51;
    ram_cell[     684] = 32'h00b89a2f;
    ram_cell[     685] = 32'h6ac68dcb;
    ram_cell[     686] = 32'h141d39a3;
    ram_cell[     687] = 32'h9d49e498;
    ram_cell[     688] = 32'h808cdf2d;
    ram_cell[     689] = 32'h256d1dee;
    ram_cell[     690] = 32'h47eab573;
    ram_cell[     691] = 32'habf5a55f;
    ram_cell[     692] = 32'h63ba2089;
    ram_cell[     693] = 32'h2ccffb64;
    ram_cell[     694] = 32'ha173712b;
    ram_cell[     695] = 32'h78c1598d;
    ram_cell[     696] = 32'he74edbe0;
    ram_cell[     697] = 32'he5886a85;
    ram_cell[     698] = 32'he26968f1;
    ram_cell[     699] = 32'h6d2b7793;
    ram_cell[     700] = 32'h72cd1f65;
    ram_cell[     701] = 32'h3eab3a5a;
    ram_cell[     702] = 32'h613f7f19;
    ram_cell[     703] = 32'hffbe8da4;
    ram_cell[     704] = 32'h7c9da6c5;
    ram_cell[     705] = 32'he2fff78b;
    ram_cell[     706] = 32'hcbdb1e4a;
    ram_cell[     707] = 32'h1ba9bdc2;
    ram_cell[     708] = 32'h55ec93ee;
    ram_cell[     709] = 32'h4058fe3e;
    ram_cell[     710] = 32'h9e3fc73b;
    ram_cell[     711] = 32'h0585eab8;
    ram_cell[     712] = 32'h4daf0c10;
    ram_cell[     713] = 32'h5e0cda18;
    ram_cell[     714] = 32'hc6a91cc4;
    ram_cell[     715] = 32'hc5efb3f7;
    ram_cell[     716] = 32'h70d39d80;
    ram_cell[     717] = 32'h7f719a12;
    ram_cell[     718] = 32'h12639c7c;
    ram_cell[     719] = 32'hc1341331;
    ram_cell[     720] = 32'h51c188fb;
    ram_cell[     721] = 32'hf847715d;
    ram_cell[     722] = 32'h1cdb5539;
    ram_cell[     723] = 32'h3274ba69;
    ram_cell[     724] = 32'h13d4fc77;
    ram_cell[     725] = 32'hed4b23c4;
    ram_cell[     726] = 32'h238c5f91;
    ram_cell[     727] = 32'h6940ad99;
    ram_cell[     728] = 32'h596f0da0;
    ram_cell[     729] = 32'h3bf1951a;
    ram_cell[     730] = 32'h29ba12ef;
    ram_cell[     731] = 32'h19af7ef3;
    ram_cell[     732] = 32'h24ecba92;
    ram_cell[     733] = 32'h80baa3b5;
    ram_cell[     734] = 32'h42808836;
    ram_cell[     735] = 32'hf3b3bd4f;
    ram_cell[     736] = 32'hecf20fc6;
    ram_cell[     737] = 32'h016765ea;
    ram_cell[     738] = 32'h13192664;
    ram_cell[     739] = 32'hcc778da9;
    ram_cell[     740] = 32'h93257bc0;
    ram_cell[     741] = 32'h006ad1c5;
    ram_cell[     742] = 32'h4a096e17;
    ram_cell[     743] = 32'hb9c7f42d;
    ram_cell[     744] = 32'h2bea556d;
    ram_cell[     745] = 32'h51083974;
    ram_cell[     746] = 32'hff3183bc;
    ram_cell[     747] = 32'h9923576e;
    ram_cell[     748] = 32'h851b7e06;
    ram_cell[     749] = 32'hf45df914;
    ram_cell[     750] = 32'h1e05b6f9;
    ram_cell[     751] = 32'h0cb1ffd2;
    ram_cell[     752] = 32'hd9bb88ff;
    ram_cell[     753] = 32'h6165d221;
    ram_cell[     754] = 32'hc5365c59;
    ram_cell[     755] = 32'hb6b02f05;
    ram_cell[     756] = 32'h09619c30;
    ram_cell[     757] = 32'h4e11cf49;
    ram_cell[     758] = 32'h83a9eae7;
    ram_cell[     759] = 32'he7078a50;
    ram_cell[     760] = 32'h4dc30d69;
    ram_cell[     761] = 32'h24a75db5;
    ram_cell[     762] = 32'ha3bb5cda;
    ram_cell[     763] = 32'h3d598231;
    ram_cell[     764] = 32'h04ed14df;
    ram_cell[     765] = 32'he937f7f9;
    ram_cell[     766] = 32'he5cc2bde;
    ram_cell[     767] = 32'h1d5fd9d0;
end

endmodule

