////////////////////////////////////////////////////////////////////////////////
// Engineer:       Jiang Binze - jiangbinze@mail.ustc.edu.cn                  //
//                                                                            //
// Design Name:    Top level module                                           //
// Project Name:   RISCV Core                                                 //
// Language:       SystemVerilog                                              //
//                                                                            //
// Description:    Top level module of the RISC-V core.                       //
//                                                                            //
////////////////////////////////////////////////////////////////////////////////

module RV32Core import core_pkg::*;
#(
    parameter DEBUG             = 1,
    parameter USE_RAM_IP        = 0,
    parameter USE_CACHE         = 1,
    parameter USE_BTB           = 1,
    parameter USE_BHT           = 0
)
(
    input   logic           clk,
    input   logic           rst,

    output  logic   [15:0]  LED

    // // Debug Signals
    // input   logic   [31:0]  CPU_Debug_DataRAM_A2,
    // input   logic   [31:0]  CPU_Debug_DataRAM_WD2,
    // input   logic   [3 :0]  CPU_Debug_DataRAM_WE2,
    // output  logic   [31:0]  CPU_Debug_DataRAM_RD2,
    // input   logic   [31:0]  CPU_Debug_InstRAM_A2,
    // input   logic   [31:0]  CPU_Debug_InstRAM_WD2,
    // input   logic   [3 :0]  CPU_Debug_InstRAM_WE2,
    // output  logic   [31:0]  CPU_Debug_InstRAM_RD2
);

    logic   [31:0]  pc_if;
    logic   [31:0]  pc_id;
    logic   [31:0]  pc_ex;
    logic   [31:0]  pc_me;
    // logic   [31:0]  pc_wb; // pc_wb is in WB module

    logic           stall_if;
    logic           stall_id;
    logic           stall_ex;
    logic           stall_me;
    logic           stall_wb;
    logic           clear_if;
    logic           clear_id;
    logic           clear_ex;
    logic           clear_me;
    logic           clear_wb;

    // IF-ID
    logic           branch_prediction_if;
    
    // ID-EX
    logic           alu_ex_ex;
    logic   [ALU_OP_WIDTH-1:0]  alu_op_ex;
    logic   [ALU_SRC_WIDTH-1:0] alu_src_1_ex;
    logic   [ALU_SRC_WIDTH-1:0] alu_src_2_ex;
    logic   [4 :0]  rs1_raddr_ex;
    logic   [4 :0]  rs2_raddr_ex;
    logic   [31:0]  rs1_rdata_ex;
    logic   [31:0]  rs2_rdata_ex;
    logic           rs1_used_ex;
    logic           rs2_used_ex;
    logic   [31:0]  imm_ex;
    logic   [4 :0]  regfile_waddr_ex;
    logic           regfile_we_ex;
    logic   [WB_WR_MUX_OP_WIDTH-1:0] regfile_wr_mux_ex;
    logic           mem_req_ex;
    logic           mem_we_ex;
    logic   [2 :0]  mem_type_ex;
    logic   [BRCH_OP_WIDTH-1:0] branch_type_ex;
    logic   [CSR_ADDR_WIDTH-1:0] csr_addr_ex;
    logic   [2 :0]  csr_type_ex;
    logic           csr_we_ex;
    logic           branch_predicition_ex;

    // EX-MEM
    logic   [31:0]  alu_result_mem;
    logic   [4 :0]  regfile_waddr_mem;
    logic           regfile_we_mem;
    logic   [WB_WR_MUX_OP_WIDTH-1:0] regfile_wr_mux_mem;
    logic           mem_req_mem;
    logic           mem_we_mem;
    logic   [2 :0]  mem_type_mem;
    logic   [31:0]  mem_wdata_mem;

    // MEM-WB
    logic           mem_req_wb;
    logic           mem_we_wb;
    logic   [3 :0]  mem_be_wb;
    logic   [2 :0]  mem_type_wb;
    logic   [31:0]  mem_addr_wb;
    logic   [31:0]  mem_wdata_wb;
    logic   [4 :0]  regfile_waddr_wb;
    logic   [31:0]  regfile_wdata_wb;
    logic           regfile_we_wb;
    logic   [WB_WR_MUX_OP_WIDTH-1:0] regfile_wr_mux_wb;

    // WB out
    logic   [4 :0]  regfile_waddr;
    logic   [31:0]  regfile_wdata;
    logic           regfile_we;

    // TO Controller
    logic           jump_decision;
    logic           branch_decision;
    logic           pc_set;
    logic   [3 :0]  pc_mux;
    logic   [4 :0]  rs1_raddr;
    logic   [4 :0]  rs2_raddr;
    logic           rs1_used;
    logic           rs2_used;
    logic           mem_req;
    logic   [4 :0]  regfile_waddr_ctrl_m;
    logic           regfile_we_ctrl_m;
    logic   [4 :0]  regfile_waddr_ctrl_w;
    logic           regfile_we_ctrl_w;
    logic           mem_miss;
    logic           branch_prediction;
    logic           branch_in_ex;
    logic   [BRCH_OP_WIDTH-1:0] branch_type;

    // Forward signals
    logic   [31:0]  regfile_wdata_fw_mem;
    logic   [31:0]  regfile_wdata_fw_wb;
    logic   [1 :0]  rs1_forward;
    logic   [1 :0]  rs2_forward;
    // Jumps and Branches
    logic   [31:0]  jump_target;
    logic   [31:0]  branch_target;
    // BTB and BHT 
    // logic   [31:0]  btb_pc_brancher;
    logic           btb_pc_we;
    // logic   [31:0]  btb_pc_target;
    logic           btb_pc_clear;
    // logic   [31:0]  bht_pc_brancher;
    logic           bht_branch_prediction;
    logic           bht_we;

    assign regfile_wdata_fw_wb  = regfile_wdata;
    assign regfile_waddr_ctrl_w = regfile_waddr;
    assign regfile_we_ctrl_w    = regfile_we;

    assign LED = pc_if[15:0];

  //////////////////////////////////////////////////
  //   ___ _____   ____ _____  _    ____ _____    //
  //  |_ _|  ___| / ___|_   _|/ \  / ___| ____|   //
  //   | || |_    \___ \ | | / _ \| |  _|  _|     //
  //   | ||  _|    ___) || |/ ___ \ |_| | |___    //
  //  |___|_|     |____/ |_/_/   \_\____|_____|   //
  //                                              //
  //////////////////////////////////////////////////
    if_stage
    #(
        .DEBUG              ( DEBUG             ),
        .USE_BTB            ( USE_BTB           ),
        .USE_BHT            ( USE_BHT           )
    )
    if_stage_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),

        .stall_if_i         ( stall_if          ),
        .clear_if_i         ( clear_if          ),

        .pc_set_i           ( pc_set            ),
        .pc_mux_i           ( pc_mux            ),
        .pc_ex_i            ( pc_ex             ),
        .boot_addr_i        ( 32'h0             ),
        .jump_target_id_i   ( jump_target       ),
        .branch_target_ex_i ( branch_target     ),

        // IF-ID Pipeline
        .pc_if_o            ( pc_if             ),
        .branch_prediction_if_o(branch_prediction_if),
        
        // branch prediction wires
        .btb_pc_brancher_i  ( pc_ex             ),
        .btb_pc_we_i        ( btb_pc_we         ),
        .btb_pc_target_i    ( branch_target     ),
        .btb_pc_clear_i     ( btb_pc_clear      ),

        .bht_pc_brancher_i  ( pc_ex             ),
        .bht_branch_deicision_i(bht_branch_prediction),
        .bht_we_i           ( bht_we            )
    ); 

  /////////////////////////////////////////////////
  //   ___ ____    ____ _____  _    ____ _____   //
  //  |_ _|  _ \  / ___|_   _|/ \  / ___| ____|  //
  //   | || | | | \___ \ | | / _ \| |  _|  _|    //
  //   | || |_| |  ___) || |/ ___ \ |_| | |___   //
  //  |___|____/  |____/ |_/_/   \_\____|_____|  //
  //                                             //
  /////////////////////////////////////////////////
    id_stage
    #(
        .DEBUG              ( DEBUG             ),
        .USE_RAM_IP         ( USE_RAM_IP        ),
        .USE_CACHE          ( USE_CACHE         ),
        .USE_BTB            ( USE_BTB           ),
        .USE_BHT            ( USE_BHT           )

    )
    id_stage_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),

        .stall_id_i         ( stall_id          ),
        .clear_id_i         ( clear_id          ),

        // From IF stage
        .pc_if_i            ( pc_if             ),
        .branch_prediction_if_i(branch_prediction_if),

        // jumps in id
        .jump_decision_o    ( jump_decision     ),
        .jump_target_o      ( jump_target       ),

        // ID-EX Pipeline
        .pc_id_o            ( pc_id             ),
        .alu_en_ex_o        ( alu_en_ex         ),
        .alu_op_ex_o        ( alu_op_ex         ),
        .alu_src_1_ex_o     ( alu_src_1_ex      ),
        .alu_src_2_ex_o     ( alu_src_2_ex      ),
        .rs1_raddr_ex_o     ( rs1_raddr_ex      ),
        .rs2_raddr_ex_o     ( rs2_raddr_ex      ),
        .rs1_rdata_ex_o     ( rs1_rdata_ex      ),
        .rs2_rdata_ex_o     ( rs2_rdata_ex      ),
        .rs1_used_ex_o      ( rs1_used_ex       ),
        .rs2_used_ex_o      ( rs2_used_ex       ),
        .imm_ex_o           ( imm_ex            ),
        .regfile_waddr_ex_o ( regfile_waddr_ex  ),
        .regfile_we_ex_o    ( regfile_we_ex     ),
        .regfile_wr_mux_ex_o( regfile_wr_mux_ex ),
        .mem_req_ex_o       ( mem_req_ex        ),
        .mem_we_ex_o        ( mem_we_ex         ),
        .mem_type_ex_o      ( mem_type_ex       ),
        .branch_type_ex_o   ( branch_type_ex    ),
        .csr_addr_ex_o      ( csr_addr_ex       ),
        .csr_we_ex_o        ( csr_we_ex         ),
        .csr_type_ex_o      ( csr_type_ex       ),
        .branch_prediction_ex_o(branch_prediction_ex),

        // From WB stage
        .regfile_waddr_wb_i ( regfile_waddr     ),
        .regfile_we_wb_i    ( regfile_we        ),
        .regfile_wdata_wb_i ( regfile_wdata     )
    );

  /////////////////////////////////////////////////////
  //   _______  __  ____ _____  _    ____ _____      //
  //  | ____\ \/ / / ___|_   _|/ \  / ___| ____|     //
  //  |  _|  \  /  \___ \ | | / _ \| |  _|  _|       //
  //  | |___ /  \   ___) || |/ ___ \ |_| | |___      //
  //  |_____/_/\_\ |____/ |_/_/   \_\____|_____|     //
  //                                                 //
  /////////////////////////////////////////////////////
    ex_stage
    #(
        .DEBUG              ( DEBUG             ),
        .USE_BTB            ( USE_BTB           ),
        .USE_BHT            ( USE_BHT           )

    )
    ex_stage_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),

        .stall_ex_i         ( stall_ex          ),
        .clear_ex_i         ( clear_ex          ),

        // From ID stage
        .pc_id_i            ( pc_id             ),
        .alu_en_i           ( alu_en_ex         ),       
        .alu_op_i           ( alu_op_ex         ),
        .alu_src_1_i        ( alu_src_1_ex      ),
        .alu_src_2_i        ( alu_src_2_ex      ),
        .rs1_raddr_i        ( rs1_raddr_ex      ),
        .rs2_raddr_i        ( rs2_raddr_ex      ),
        .rs1_rdata_i        ( rs1_rdata_ex      ),
        .rs2_rdata_i        ( rs2_rdata_ex      ),
        .rs1_used_i         ( rs1_used_ex       ),
        .rs2_used_i         ( rs2_used_ex       ),
        .imm_i              ( imm_ex            ),
        .regfile_waddr_i    ( regfile_waddr_ex  ),
        .regfile_we_i       ( regfile_we_ex     ),
        .regfile_wr_mux_i   ( regfile_wr_mux_ex ),
        .mem_req_i          ( mem_req_ex        ),
        .mem_we_i           ( mem_we_ex         ),
        .mem_type_i         ( mem_type_ex       ),
        .branch_type_i      ( branch_type_ex    ),
        .csr_addr_i         ( csr_addr_ex       ),
        .csr_type_i         ( csr_type_ex       ),
        .csr_we_i           ( csr_we_ex         ),
        .branch_prediction_i(branch_prediction_ex),

        // handle branches
        .branch_decision_o  ( branch_decision   ),
        .branch_target_o    ( branch_target     ),
        .branch_prediction_o( branch_prediction ),
        .branch_in_ex_o     ( branch_in_ex      ),
        .branch_type_o      ( branch_type       ),

        // to controller
        .rs1_raddr_o        ( rs1_raddr         ),
        .rs2_raddr_o        ( rs2_raddr         ),
        .rs1_used_o         ( rs1_used          ),
        .rs2_used_o         ( rs2_used          ),

        // EX-MEM Pipeline
        .pc_ex_o            ( pc_ex             ),
        .alu_result_mem_o   ( alu_result_mem    ),
        .regfile_waddr_mem_o( regfile_waddr_mem ),
        .regfile_we_mem_o   ( regfile_we_mem    ),
        .regfile_wr_mux_mem_o(regfile_wr_mux_mem),
        .mem_req_mem_o      ( mem_req_mem       ),
        .mem_we_mem_o       ( mem_we_mem        ),
        .mem_type_mem_o     ( mem_type_mem      ),
        .mem_wdata_mem_o    ( mem_wdata_mem     ),
        
        // Forward Data
        .regfile_wdata_mem_i( regfile_wdata_fw_mem),
        .regfile_wdata_wb_i ( regfile_wdata_fw_wb ),
        .rs1_forward_i      ( rs1_forward       ),
        .rs2_forward_i      ( rs2_forward       )
    );

    // MEM stage
    mem_stage
    #( 
        .DEBUG              ( DEBUG             )
    )
    mem_stage_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),

        .stall_mem_i        ( stall_me          ),
        .clear_mem_i        ( clear_me          ),

        // From EX
        .pc_ex_i            ( pc_ex             ),
        .alu_result_i       ( alu_result_mem    ),
        .regfile_waddr_i    ( regfile_waddr_mem ),
        .regfile_we_i       ( regfile_we_mem    ),
        .regfile_wr_mux_i   ( regfile_wr_mux_mem),
        .mem_req_i          ( mem_req_mem       ),
        .mem_we_i           ( mem_we_mem        ),
        .mem_type_i         ( mem_type_mem      ),
        .mem_wdata_i        ( mem_wdata_mem     ),

        // to controller
        .mem_req_o          ( mem_req           ),    // used to justify whether it is a load instr
        .regfile_waddr_o    ( regfile_waddr_ctrl_m),
        .regfile_we_o       ( regfile_we_ctrl_m),
        // forward
        .regfile_wdata_o    ( regfile_wdata_fw_mem),

        // MEM-WB Pipeline
        .pc_mem_o           ( pc_me             ),
        .mem_req_wb_o       ( mem_req_wb        ), 
        .mem_we_wb_o        ( mem_we_wb         ),
        .mem_be_wb_o        ( mem_be_wb         ),
        .mem_type_wb_o      ( mem_type_wb       ),
        .mem_addr_wb_o      ( mem_addr_wb       ),
        .mem_wdata_wb_o     ( mem_wdata_wb      ),
        .regfile_waddr_wb_o ( regfile_waddr_wb  ),
        .regfile_wdata_wb_o ( regfile_wdata_wb  ),
        .regfile_we_wb_o    ( regfile_we_wb     ),
        .regfile_wr_mux_wb_o( regfile_wr_mux_wb )
    );

    // WB stage
    wb_stage
    #(
        .DEBUG              ( DEBUG             ),
        .USE_RAM_IP         ( USE_RAM_IP        ),
        .USE_CACHE          ( USE_CACHE         )
    )
    wb_stage_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),
        
        .stall_wb_i         ( stall_wb          ),
        .clear_wb_i         ( clear_wb          ),

        // From MEM
        .pc_mem_i           ( pc_me             ),
        .mem_req_i          ( mem_req_wb        ),
        .mem_we_i           ( mem_we_wb         ),
        .mem_be_i           ( mem_be_wb         ),
        .mem_type_i         ( mem_type_wb       ),
        .mem_addr_i         ( mem_addr_wb       ),
        .mem_wdata_i        ( mem_wdata_wb      ),
        .regfile_waddr_i    ( regfile_waddr_wb  ),
        .regfile_wdata_i    ( regfile_wdata_wb  ),
        .regfile_we_i       ( regfile_we_wb     ),
        .regfile_wr_mux_i   ( regfile_wr_mux_wb ),

        // out
        .regfile_waddr_o    ( regfile_waddr     ),
        .regfile_wdata_o    ( regfile_wdata     ),
        .regfile_we_o       ( regfile_we        ),

        .miss               ( mem_miss          )
    );

  ////////////////////////////////////////////////////////////////////
  //    ____ ___  _   _ _____ ____   ___  _     _     _____ ____    //
  //   / ___/ _ \| \ | |_   _|  _ \ / _ \| |   | |   | ____|  _ \   //
  //  | |  | | | |  \| | | | | |_) | | | | |   | |   |  _| | |_) |  //
  //  | |__| |_| | |\  | | | |  _ <| |_| | |___| |___| |___|  _ <   //
  //   \____\___/|_| \_| |_| |_| \_\\___/|_____|_____|_____|_| \_\  //
  //                                                                //
  ////////////////////////////////////////////////////////////////////
    controller 
    #(
        .DEBUG              ( DEBUG             ),
        .USE_BTB            ( USE_BTB           ),
        .USE_BHT            ( USE_BHT           )
    )
    controller_i
    (
        .clk                ( clk           ),
        .rst_n              ( ~rst          ),

        // branches and jumps
        .jump_decision_i    ( jump_decision     ),
        .branch_decision_i  ( branch_decision   ),
        .branch_prediction_i( branch_prediction ),
        .branch_in_ex_i     ( branch_in_ex      ),
        .branch_type_i      ( branch_type       ),
        .pc_set_o           ( pc_set            ),
        .pc_mux_o           ( pc_mux            ),
        // branch_predictions
        .btb_pc_we_o        ( btb_pc_we         ),
        .btb_pc_clear_o     ( btb_pc_clear      ),
        .bht_branch_prediction_o(bht_branch_prediction),
        .bht_we_o           ( bht_we            ),

        // pipeline stall, clear signals
        .stall_if_o         ( stall_if          ),
        .stall_id_o         ( stall_id          ),
        .stall_ex_o         ( stall_ex          ),
        .stall_mem_o        ( stall_me          ),
        .stall_wb_o         ( stall_wb          ),
        .clear_if_o         ( clear_if          ),
        .clear_id_o         ( clear_id          ),
        .clear_ex_o         ( clear_ex          ),
        .clear_mem_o        ( clear_me          ),
        .clear_wb_o         ( clear_wb          ),

        // ex, mem, wb info
        .rs1_raddr_ex_i     ( rs1_raddr         ),
        .rs2_raddr_ex_i     ( rs2_raddr         ),
        .rs1_used_ex_i      ( rs1_used          ),
        .rs2_used_ex_i      ( rs2_used          ),
        .mem_req_i          ( mem_req           ),
        .regfile_waddr_mem_i( regfile_waddr_ctrl_m),
        .regfile_we_mem_i   ( regfile_we_ctrl_m),
        .regfile_waddr_wb_i ( regfile_waddr_ctrl_w),
        .regfile_we_wb_i    ( regfile_we_ctrl_w),

        // forward signals
        .rs1_forward_o      ( rs1_forward       ),
        .rs2_forward_o      ( rs2_forward       ),

        .mem_miss_i         ( mem_miss          )
    );

endmodule
