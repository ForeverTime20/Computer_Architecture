
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h9e0e9c03;
    ram_cell[       1] = 32'h0;  // 32'hc2069c70;
    ram_cell[       2] = 32'h0;  // 32'h4337cd6e;
    ram_cell[       3] = 32'h0;  // 32'h7c4af4a2;
    ram_cell[       4] = 32'h0;  // 32'hb7bb79cc;
    ram_cell[       5] = 32'h0;  // 32'h879a3d1e;
    ram_cell[       6] = 32'h0;  // 32'hf4d7feb1;
    ram_cell[       7] = 32'h0;  // 32'hecc7e06f;
    ram_cell[       8] = 32'h0;  // 32'h8c324064;
    ram_cell[       9] = 32'h0;  // 32'hd4f1ac4f;
    ram_cell[      10] = 32'h0;  // 32'h7a7bf755;
    ram_cell[      11] = 32'h0;  // 32'h3b72a8b1;
    ram_cell[      12] = 32'h0;  // 32'hb3eea433;
    ram_cell[      13] = 32'h0;  // 32'h7f4e6a4c;
    ram_cell[      14] = 32'h0;  // 32'ha3a03c26;
    ram_cell[      15] = 32'h0;  // 32'h14f27b72;
    ram_cell[      16] = 32'h0;  // 32'ha4c8af88;
    ram_cell[      17] = 32'h0;  // 32'hafea9ada;
    ram_cell[      18] = 32'h0;  // 32'hd01c60f0;
    ram_cell[      19] = 32'h0;  // 32'h46ebf5e3;
    ram_cell[      20] = 32'h0;  // 32'h9f6756e9;
    ram_cell[      21] = 32'h0;  // 32'h4e98fa08;
    ram_cell[      22] = 32'h0;  // 32'hd6d17c80;
    ram_cell[      23] = 32'h0;  // 32'hefb68c87;
    ram_cell[      24] = 32'h0;  // 32'h2cfddbb2;
    ram_cell[      25] = 32'h0;  // 32'h4ae16f17;
    ram_cell[      26] = 32'h0;  // 32'h52f8693e;
    ram_cell[      27] = 32'h0;  // 32'h7f2f19b1;
    ram_cell[      28] = 32'h0;  // 32'h148f1053;
    ram_cell[      29] = 32'h0;  // 32'h2bada337;
    ram_cell[      30] = 32'h0;  // 32'h1e865cb4;
    ram_cell[      31] = 32'h0;  // 32'hc41e2614;
    ram_cell[      32] = 32'h0;  // 32'h722779a1;
    ram_cell[      33] = 32'h0;  // 32'hea9e2198;
    ram_cell[      34] = 32'h0;  // 32'h63002d5b;
    ram_cell[      35] = 32'h0;  // 32'h37d99548;
    ram_cell[      36] = 32'h0;  // 32'ha24dbf88;
    ram_cell[      37] = 32'h0;  // 32'h8fc20020;
    ram_cell[      38] = 32'h0;  // 32'h7b920ddd;
    ram_cell[      39] = 32'h0;  // 32'h10198b6e;
    ram_cell[      40] = 32'h0;  // 32'h0198ce7d;
    ram_cell[      41] = 32'h0;  // 32'h8d6ccdaa;
    ram_cell[      42] = 32'h0;  // 32'hd412a7a0;
    ram_cell[      43] = 32'h0;  // 32'hc35a6e2d;
    ram_cell[      44] = 32'h0;  // 32'hcd338b48;
    ram_cell[      45] = 32'h0;  // 32'h2bbcbb2b;
    ram_cell[      46] = 32'h0;  // 32'hcedf7b70;
    ram_cell[      47] = 32'h0;  // 32'h544fc389;
    ram_cell[      48] = 32'h0;  // 32'h8160b4b6;
    ram_cell[      49] = 32'h0;  // 32'h61470c3b;
    ram_cell[      50] = 32'h0;  // 32'hf58bddbe;
    ram_cell[      51] = 32'h0;  // 32'h24b76488;
    ram_cell[      52] = 32'h0;  // 32'h1eba8020;
    ram_cell[      53] = 32'h0;  // 32'h3e70db0f;
    ram_cell[      54] = 32'h0;  // 32'h18ef112b;
    ram_cell[      55] = 32'h0;  // 32'h2f51ecaa;
    ram_cell[      56] = 32'h0;  // 32'ha17196f5;
    ram_cell[      57] = 32'h0;  // 32'h8938888c;
    ram_cell[      58] = 32'h0;  // 32'h33b9bbdc;
    ram_cell[      59] = 32'h0;  // 32'he5efe63d;
    ram_cell[      60] = 32'h0;  // 32'h0a61cdf0;
    ram_cell[      61] = 32'h0;  // 32'h091b8fbe;
    ram_cell[      62] = 32'h0;  // 32'h7c1a1283;
    ram_cell[      63] = 32'h0;  // 32'h7e505d38;
    ram_cell[      64] = 32'h0;  // 32'h58f01d01;
    ram_cell[      65] = 32'h0;  // 32'h78066e85;
    ram_cell[      66] = 32'h0;  // 32'hddee3c98;
    ram_cell[      67] = 32'h0;  // 32'h39ad7ca5;
    ram_cell[      68] = 32'h0;  // 32'hb04cfea6;
    ram_cell[      69] = 32'h0;  // 32'hba4416fb;
    ram_cell[      70] = 32'h0;  // 32'h095907a9;
    ram_cell[      71] = 32'h0;  // 32'h8e59d1d7;
    ram_cell[      72] = 32'h0;  // 32'hc1522a06;
    ram_cell[      73] = 32'h0;  // 32'h1e7934fa;
    ram_cell[      74] = 32'h0;  // 32'h4636e20d;
    ram_cell[      75] = 32'h0;  // 32'h12860053;
    ram_cell[      76] = 32'h0;  // 32'h9233fbaa;
    ram_cell[      77] = 32'h0;  // 32'h4e1b695a;
    ram_cell[      78] = 32'h0;  // 32'h8c22e8e4;
    ram_cell[      79] = 32'h0;  // 32'h47d317f5;
    ram_cell[      80] = 32'h0;  // 32'hb6d3a71c;
    ram_cell[      81] = 32'h0;  // 32'h86a98f2b;
    ram_cell[      82] = 32'h0;  // 32'h3e09fcd3;
    ram_cell[      83] = 32'h0;  // 32'hbf1deb92;
    ram_cell[      84] = 32'h0;  // 32'hf693a0e5;
    ram_cell[      85] = 32'h0;  // 32'hb664b924;
    ram_cell[      86] = 32'h0;  // 32'h96445315;
    ram_cell[      87] = 32'h0;  // 32'h41ae867e;
    ram_cell[      88] = 32'h0;  // 32'h937177b2;
    ram_cell[      89] = 32'h0;  // 32'h56387ba2;
    ram_cell[      90] = 32'h0;  // 32'h2d5a0873;
    ram_cell[      91] = 32'h0;  // 32'he1843c36;
    ram_cell[      92] = 32'h0;  // 32'hb546fdac;
    ram_cell[      93] = 32'h0;  // 32'hf2cbc11f;
    ram_cell[      94] = 32'h0;  // 32'h2a49eadc;
    ram_cell[      95] = 32'h0;  // 32'h09aad16c;
    ram_cell[      96] = 32'h0;  // 32'h932e833d;
    ram_cell[      97] = 32'h0;  // 32'h65ff55a9;
    ram_cell[      98] = 32'h0;  // 32'hb1977045;
    ram_cell[      99] = 32'h0;  // 32'h72038cce;
    ram_cell[     100] = 32'h0;  // 32'h0444b59f;
    ram_cell[     101] = 32'h0;  // 32'h05e7f528;
    ram_cell[     102] = 32'h0;  // 32'h153f38a1;
    ram_cell[     103] = 32'h0;  // 32'h071fd09b;
    ram_cell[     104] = 32'h0;  // 32'hf40a1202;
    ram_cell[     105] = 32'h0;  // 32'h22056c95;
    ram_cell[     106] = 32'h0;  // 32'h17655632;
    ram_cell[     107] = 32'h0;  // 32'h5b76152a;
    ram_cell[     108] = 32'h0;  // 32'h107e2084;
    ram_cell[     109] = 32'h0;  // 32'h4a75aaf0;
    ram_cell[     110] = 32'h0;  // 32'hf6999682;
    ram_cell[     111] = 32'h0;  // 32'h59ed10f4;
    ram_cell[     112] = 32'h0;  // 32'hb9380597;
    ram_cell[     113] = 32'h0;  // 32'h1d96dadf;
    ram_cell[     114] = 32'h0;  // 32'h9e0f44cd;
    ram_cell[     115] = 32'h0;  // 32'h904010d9;
    ram_cell[     116] = 32'h0;  // 32'hb4c82ab8;
    ram_cell[     117] = 32'h0;  // 32'h5bcdb8b2;
    ram_cell[     118] = 32'h0;  // 32'h0856fa5a;
    ram_cell[     119] = 32'h0;  // 32'h8b0a52b7;
    ram_cell[     120] = 32'h0;  // 32'h62507cf8;
    ram_cell[     121] = 32'h0;  // 32'hf361bac6;
    ram_cell[     122] = 32'h0;  // 32'h3b27b530;
    ram_cell[     123] = 32'h0;  // 32'h2ef26d1a;
    ram_cell[     124] = 32'h0;  // 32'he863bfb8;
    ram_cell[     125] = 32'h0;  // 32'h1eebea54;
    ram_cell[     126] = 32'h0;  // 32'hac60f04a;
    ram_cell[     127] = 32'h0;  // 32'h14553e53;
    ram_cell[     128] = 32'h0;  // 32'ha3c82f1a;
    ram_cell[     129] = 32'h0;  // 32'hfc6014f6;
    ram_cell[     130] = 32'h0;  // 32'h63c5ac0e;
    ram_cell[     131] = 32'h0;  // 32'h039e819f;
    ram_cell[     132] = 32'h0;  // 32'hf8658187;
    ram_cell[     133] = 32'h0;  // 32'hb0191252;
    ram_cell[     134] = 32'h0;  // 32'h701f9bdf;
    ram_cell[     135] = 32'h0;  // 32'h41065223;
    ram_cell[     136] = 32'h0;  // 32'hbd9cfc60;
    ram_cell[     137] = 32'h0;  // 32'hb54c5bce;
    ram_cell[     138] = 32'h0;  // 32'hfb8e4ec3;
    ram_cell[     139] = 32'h0;  // 32'h24b6a65d;
    ram_cell[     140] = 32'h0;  // 32'hc58595e6;
    ram_cell[     141] = 32'h0;  // 32'ha68847cd;
    ram_cell[     142] = 32'h0;  // 32'h9b81dd41;
    ram_cell[     143] = 32'h0;  // 32'h74e5cdb2;
    ram_cell[     144] = 32'h0;  // 32'h63932a79;
    ram_cell[     145] = 32'h0;  // 32'h1bc7fccc;
    ram_cell[     146] = 32'h0;  // 32'h6daad863;
    ram_cell[     147] = 32'h0;  // 32'h294989f6;
    ram_cell[     148] = 32'h0;  // 32'h23a4fd4c;
    ram_cell[     149] = 32'h0;  // 32'h42d9e5d8;
    ram_cell[     150] = 32'h0;  // 32'h319bc775;
    ram_cell[     151] = 32'h0;  // 32'h7dec53e9;
    ram_cell[     152] = 32'h0;  // 32'h46fab970;
    ram_cell[     153] = 32'h0;  // 32'he6529b3a;
    ram_cell[     154] = 32'h0;  // 32'h675ce968;
    ram_cell[     155] = 32'h0;  // 32'h5c0a13df;
    ram_cell[     156] = 32'h0;  // 32'h5d9ab324;
    ram_cell[     157] = 32'h0;  // 32'h41166e71;
    ram_cell[     158] = 32'h0;  // 32'h5bd0baed;
    ram_cell[     159] = 32'h0;  // 32'h5af7bbfd;
    ram_cell[     160] = 32'h0;  // 32'h2d273a64;
    ram_cell[     161] = 32'h0;  // 32'h3e49bb70;
    ram_cell[     162] = 32'h0;  // 32'hd10788ad;
    ram_cell[     163] = 32'h0;  // 32'h526b4517;
    ram_cell[     164] = 32'h0;  // 32'h86048562;
    ram_cell[     165] = 32'h0;  // 32'h90a3fa7d;
    ram_cell[     166] = 32'h0;  // 32'hc76c6fe0;
    ram_cell[     167] = 32'h0;  // 32'h130bb17e;
    ram_cell[     168] = 32'h0;  // 32'h34281913;
    ram_cell[     169] = 32'h0;  // 32'h238bb28f;
    ram_cell[     170] = 32'h0;  // 32'h3ceb4d69;
    ram_cell[     171] = 32'h0;  // 32'he17efc65;
    ram_cell[     172] = 32'h0;  // 32'h079d13c4;
    ram_cell[     173] = 32'h0;  // 32'h7e2dcf89;
    ram_cell[     174] = 32'h0;  // 32'hb9d2c125;
    ram_cell[     175] = 32'h0;  // 32'h4992409d;
    ram_cell[     176] = 32'h0;  // 32'h9ec5ac31;
    ram_cell[     177] = 32'h0;  // 32'h57fb3816;
    ram_cell[     178] = 32'h0;  // 32'hcd136ce1;
    ram_cell[     179] = 32'h0;  // 32'h3307b7dd;
    ram_cell[     180] = 32'h0;  // 32'h68a09a41;
    ram_cell[     181] = 32'h0;  // 32'hd7bf5f69;
    ram_cell[     182] = 32'h0;  // 32'h422c2d64;
    ram_cell[     183] = 32'h0;  // 32'h2750b435;
    ram_cell[     184] = 32'h0;  // 32'h23a59ec5;
    ram_cell[     185] = 32'h0;  // 32'h94f40b82;
    ram_cell[     186] = 32'h0;  // 32'h4ffc5d49;
    ram_cell[     187] = 32'h0;  // 32'h22987ff9;
    ram_cell[     188] = 32'h0;  // 32'heeeaba55;
    ram_cell[     189] = 32'h0;  // 32'h05cc645a;
    ram_cell[     190] = 32'h0;  // 32'h0e3ce922;
    ram_cell[     191] = 32'h0;  // 32'hfc51a00d;
    ram_cell[     192] = 32'h0;  // 32'hafdb2747;
    ram_cell[     193] = 32'h0;  // 32'h36d9b10f;
    ram_cell[     194] = 32'h0;  // 32'hb31fbb69;
    ram_cell[     195] = 32'h0;  // 32'he04a2eec;
    ram_cell[     196] = 32'h0;  // 32'heb2edcd0;
    ram_cell[     197] = 32'h0;  // 32'hbcd2ef65;
    ram_cell[     198] = 32'h0;  // 32'hd82c624b;
    ram_cell[     199] = 32'h0;  // 32'hc2cf8e1c;
    ram_cell[     200] = 32'h0;  // 32'h50fca10e;
    ram_cell[     201] = 32'h0;  // 32'h6d2a99c6;
    ram_cell[     202] = 32'h0;  // 32'hb9d44441;
    ram_cell[     203] = 32'h0;  // 32'hca8e36c2;
    ram_cell[     204] = 32'h0;  // 32'hfc2cb380;
    ram_cell[     205] = 32'h0;  // 32'h515ecfff;
    ram_cell[     206] = 32'h0;  // 32'h3431a6bd;
    ram_cell[     207] = 32'h0;  // 32'h7fff93e1;
    ram_cell[     208] = 32'h0;  // 32'h64ac9ee1;
    ram_cell[     209] = 32'h0;  // 32'h49d69fe5;
    ram_cell[     210] = 32'h0;  // 32'hc1a01fe3;
    ram_cell[     211] = 32'h0;  // 32'h8fb31b13;
    ram_cell[     212] = 32'h0;  // 32'he99d3ef8;
    ram_cell[     213] = 32'h0;  // 32'h8ebe69d1;
    ram_cell[     214] = 32'h0;  // 32'h0fda63df;
    ram_cell[     215] = 32'h0;  // 32'h743fa243;
    ram_cell[     216] = 32'h0;  // 32'hd68b0c82;
    ram_cell[     217] = 32'h0;  // 32'h383b888f;
    ram_cell[     218] = 32'h0;  // 32'h735598d6;
    ram_cell[     219] = 32'h0;  // 32'h6765df77;
    ram_cell[     220] = 32'h0;  // 32'h56c31fdb;
    ram_cell[     221] = 32'h0;  // 32'h13dd4d04;
    ram_cell[     222] = 32'h0;  // 32'hce4f0dff;
    ram_cell[     223] = 32'h0;  // 32'hf713260a;
    ram_cell[     224] = 32'h0;  // 32'hd1863389;
    ram_cell[     225] = 32'h0;  // 32'h766e85eb;
    ram_cell[     226] = 32'h0;  // 32'hecd1dd67;
    ram_cell[     227] = 32'h0;  // 32'hbdd92016;
    ram_cell[     228] = 32'h0;  // 32'h9e8ecc00;
    ram_cell[     229] = 32'h0;  // 32'h6f7a4c80;
    ram_cell[     230] = 32'h0;  // 32'h18518fb5;
    ram_cell[     231] = 32'h0;  // 32'hdf59fdd8;
    ram_cell[     232] = 32'h0;  // 32'h88fa48ae;
    ram_cell[     233] = 32'h0;  // 32'h87aea642;
    ram_cell[     234] = 32'h0;  // 32'hb05a7794;
    ram_cell[     235] = 32'h0;  // 32'h47adfc03;
    ram_cell[     236] = 32'h0;  // 32'h2c9ccd70;
    ram_cell[     237] = 32'h0;  // 32'hc9020557;
    ram_cell[     238] = 32'h0;  // 32'h8e12f0f4;
    ram_cell[     239] = 32'h0;  // 32'h04df2b34;
    ram_cell[     240] = 32'h0;  // 32'h148e9919;
    ram_cell[     241] = 32'h0;  // 32'h39903ebc;
    ram_cell[     242] = 32'h0;  // 32'h3978789b;
    ram_cell[     243] = 32'h0;  // 32'h3d81d269;
    ram_cell[     244] = 32'h0;  // 32'h0a64786d;
    ram_cell[     245] = 32'h0;  // 32'h93e31add;
    ram_cell[     246] = 32'h0;  // 32'h678849b1;
    ram_cell[     247] = 32'h0;  // 32'hc3913752;
    ram_cell[     248] = 32'h0;  // 32'h68ccf07e;
    ram_cell[     249] = 32'h0;  // 32'h2b850be9;
    ram_cell[     250] = 32'h0;  // 32'h7f1f170f;
    ram_cell[     251] = 32'h0;  // 32'hc105dc37;
    ram_cell[     252] = 32'h0;  // 32'h135443be;
    ram_cell[     253] = 32'h0;  // 32'h69a88ed2;
    ram_cell[     254] = 32'h0;  // 32'hed3e8c7a;
    ram_cell[     255] = 32'h0;  // 32'hbe397583;
    // src matrix A
    ram_cell[     256] = 32'hdc1bf809;
    ram_cell[     257] = 32'hd8c4b5a4;
    ram_cell[     258] = 32'hf8e9eb9e;
    ram_cell[     259] = 32'haedd147f;
    ram_cell[     260] = 32'h9dac5737;
    ram_cell[     261] = 32'hcfe547d7;
    ram_cell[     262] = 32'hb6ef258c;
    ram_cell[     263] = 32'h0cdfe75b;
    ram_cell[     264] = 32'hf92c7437;
    ram_cell[     265] = 32'h16a23307;
    ram_cell[     266] = 32'h15cf4959;
    ram_cell[     267] = 32'hdd8e63f3;
    ram_cell[     268] = 32'hfbc7d95b;
    ram_cell[     269] = 32'h1b7c51e8;
    ram_cell[     270] = 32'haee0b756;
    ram_cell[     271] = 32'h250d7ae6;
    ram_cell[     272] = 32'h747d81a3;
    ram_cell[     273] = 32'h94f4b6e6;
    ram_cell[     274] = 32'h1538cf47;
    ram_cell[     275] = 32'h267bc2bb;
    ram_cell[     276] = 32'h3bf9a1b4;
    ram_cell[     277] = 32'h74ac024c;
    ram_cell[     278] = 32'h4091db28;
    ram_cell[     279] = 32'h4dc2048a;
    ram_cell[     280] = 32'h19acae12;
    ram_cell[     281] = 32'hbc9b4720;
    ram_cell[     282] = 32'hbbd0b5dc;
    ram_cell[     283] = 32'h20dc50a5;
    ram_cell[     284] = 32'h5304172e;
    ram_cell[     285] = 32'h7bde68be;
    ram_cell[     286] = 32'h6d0e9817;
    ram_cell[     287] = 32'h86837865;
    ram_cell[     288] = 32'h28c13f93;
    ram_cell[     289] = 32'ha3e49854;
    ram_cell[     290] = 32'h1ddcfdc8;
    ram_cell[     291] = 32'hbaea68aa;
    ram_cell[     292] = 32'hf1305720;
    ram_cell[     293] = 32'h442b75f8;
    ram_cell[     294] = 32'h2e3b942c;
    ram_cell[     295] = 32'h2985e9c8;
    ram_cell[     296] = 32'h872e55bc;
    ram_cell[     297] = 32'hfce8d668;
    ram_cell[     298] = 32'hc002f4f2;
    ram_cell[     299] = 32'h2f76f9bc;
    ram_cell[     300] = 32'h888e1f49;
    ram_cell[     301] = 32'h7494b9df;
    ram_cell[     302] = 32'h07bb34f8;
    ram_cell[     303] = 32'h35a776e2;
    ram_cell[     304] = 32'h02501b26;
    ram_cell[     305] = 32'hff7e23e2;
    ram_cell[     306] = 32'heefd4e8c;
    ram_cell[     307] = 32'h940b4761;
    ram_cell[     308] = 32'h0e7e8358;
    ram_cell[     309] = 32'h17d91177;
    ram_cell[     310] = 32'he7f0f97f;
    ram_cell[     311] = 32'h74eb1d24;
    ram_cell[     312] = 32'h38cef189;
    ram_cell[     313] = 32'h5ccbcae1;
    ram_cell[     314] = 32'h12497652;
    ram_cell[     315] = 32'h76b33485;
    ram_cell[     316] = 32'h624f9aed;
    ram_cell[     317] = 32'haf4a9c1e;
    ram_cell[     318] = 32'h5f320e57;
    ram_cell[     319] = 32'h58ad2f2e;
    ram_cell[     320] = 32'h4d1b58a5;
    ram_cell[     321] = 32'haf4e2470;
    ram_cell[     322] = 32'ha866215d;
    ram_cell[     323] = 32'h3cbc4ec6;
    ram_cell[     324] = 32'h237cc662;
    ram_cell[     325] = 32'hde1e7a56;
    ram_cell[     326] = 32'hc20837f1;
    ram_cell[     327] = 32'h39ffb1c6;
    ram_cell[     328] = 32'h0968b3fe;
    ram_cell[     329] = 32'hdb3a4999;
    ram_cell[     330] = 32'h2be4fad4;
    ram_cell[     331] = 32'h5c10bb68;
    ram_cell[     332] = 32'h222dcc2f;
    ram_cell[     333] = 32'h938a4b7d;
    ram_cell[     334] = 32'h2f5c9c23;
    ram_cell[     335] = 32'h4f58e845;
    ram_cell[     336] = 32'h1a5dc093;
    ram_cell[     337] = 32'h1bacd7c6;
    ram_cell[     338] = 32'h3578b5e7;
    ram_cell[     339] = 32'hdd64fcbc;
    ram_cell[     340] = 32'h0f5a0b32;
    ram_cell[     341] = 32'h2f8605ae;
    ram_cell[     342] = 32'hfde63e82;
    ram_cell[     343] = 32'h8a92d6b9;
    ram_cell[     344] = 32'hf25ac251;
    ram_cell[     345] = 32'h622f5557;
    ram_cell[     346] = 32'h429885dc;
    ram_cell[     347] = 32'h3befcfcc;
    ram_cell[     348] = 32'had33dce3;
    ram_cell[     349] = 32'h8875841a;
    ram_cell[     350] = 32'h936b5d15;
    ram_cell[     351] = 32'hff2a203d;
    ram_cell[     352] = 32'haf117c3b;
    ram_cell[     353] = 32'h3986ef52;
    ram_cell[     354] = 32'h50f36686;
    ram_cell[     355] = 32'hbceee364;
    ram_cell[     356] = 32'hcef49a36;
    ram_cell[     357] = 32'h8a2f1704;
    ram_cell[     358] = 32'h4dca8692;
    ram_cell[     359] = 32'h87576b94;
    ram_cell[     360] = 32'h0053fab8;
    ram_cell[     361] = 32'hb5a4f06d;
    ram_cell[     362] = 32'h063cef3c;
    ram_cell[     363] = 32'hce3a2e81;
    ram_cell[     364] = 32'hd4444308;
    ram_cell[     365] = 32'h3f4e2cc1;
    ram_cell[     366] = 32'h53df6206;
    ram_cell[     367] = 32'h9b1aa377;
    ram_cell[     368] = 32'h22f1b10b;
    ram_cell[     369] = 32'h1118c81c;
    ram_cell[     370] = 32'h6218b307;
    ram_cell[     371] = 32'h017f0951;
    ram_cell[     372] = 32'h35643a72;
    ram_cell[     373] = 32'h003a8760;
    ram_cell[     374] = 32'h12ca1e85;
    ram_cell[     375] = 32'h5b3311d4;
    ram_cell[     376] = 32'h1e95e489;
    ram_cell[     377] = 32'h9ac0a4f8;
    ram_cell[     378] = 32'h9defce55;
    ram_cell[     379] = 32'hd0f89b49;
    ram_cell[     380] = 32'hd779fa6f;
    ram_cell[     381] = 32'h1b7ad3d8;
    ram_cell[     382] = 32'he64e53d9;
    ram_cell[     383] = 32'h3e4d6254;
    ram_cell[     384] = 32'h4f5f0950;
    ram_cell[     385] = 32'h27074843;
    ram_cell[     386] = 32'h43b34006;
    ram_cell[     387] = 32'h8c099f8f;
    ram_cell[     388] = 32'h66010089;
    ram_cell[     389] = 32'hdfb88f54;
    ram_cell[     390] = 32'h404e4bb9;
    ram_cell[     391] = 32'h00c6606d;
    ram_cell[     392] = 32'he9a4f0f8;
    ram_cell[     393] = 32'h603eac19;
    ram_cell[     394] = 32'h27974e52;
    ram_cell[     395] = 32'he9b273c2;
    ram_cell[     396] = 32'h33293377;
    ram_cell[     397] = 32'h88ae62ad;
    ram_cell[     398] = 32'h71e7b7a3;
    ram_cell[     399] = 32'h7cc2143f;
    ram_cell[     400] = 32'hd22741c6;
    ram_cell[     401] = 32'hf436b1b6;
    ram_cell[     402] = 32'ha6f9ca1d;
    ram_cell[     403] = 32'h57e3f10d;
    ram_cell[     404] = 32'h1815eeca;
    ram_cell[     405] = 32'h3b943511;
    ram_cell[     406] = 32'hee3895cf;
    ram_cell[     407] = 32'h431f0a8d;
    ram_cell[     408] = 32'h9517b4d6;
    ram_cell[     409] = 32'h16856b37;
    ram_cell[     410] = 32'hb2e0f4e0;
    ram_cell[     411] = 32'h0da849d9;
    ram_cell[     412] = 32'h91ad21fc;
    ram_cell[     413] = 32'h1736bf3b;
    ram_cell[     414] = 32'h7e412ad0;
    ram_cell[     415] = 32'h04409ade;
    ram_cell[     416] = 32'h85c65744;
    ram_cell[     417] = 32'h3076248f;
    ram_cell[     418] = 32'h60e607c7;
    ram_cell[     419] = 32'h07956ee9;
    ram_cell[     420] = 32'hb75e947e;
    ram_cell[     421] = 32'h7348ee55;
    ram_cell[     422] = 32'h31f0bc3e;
    ram_cell[     423] = 32'h5169fcb4;
    ram_cell[     424] = 32'h85775ad2;
    ram_cell[     425] = 32'h07367ec9;
    ram_cell[     426] = 32'h95fe89a3;
    ram_cell[     427] = 32'h9f2c5f68;
    ram_cell[     428] = 32'hcf2b73a4;
    ram_cell[     429] = 32'ha7ba3aa3;
    ram_cell[     430] = 32'h40ba4849;
    ram_cell[     431] = 32'h86760386;
    ram_cell[     432] = 32'hed852820;
    ram_cell[     433] = 32'hc83a0a6b;
    ram_cell[     434] = 32'h83108472;
    ram_cell[     435] = 32'h4c2e1867;
    ram_cell[     436] = 32'h770bb2eb;
    ram_cell[     437] = 32'h97490fb8;
    ram_cell[     438] = 32'h7d0871e3;
    ram_cell[     439] = 32'h7a6bd28a;
    ram_cell[     440] = 32'h423deb51;
    ram_cell[     441] = 32'h0079f74f;
    ram_cell[     442] = 32'hd3878927;
    ram_cell[     443] = 32'h04ec6987;
    ram_cell[     444] = 32'h1b393754;
    ram_cell[     445] = 32'h3c819a4b;
    ram_cell[     446] = 32'h67441815;
    ram_cell[     447] = 32'h54a458b2;
    ram_cell[     448] = 32'h45793a14;
    ram_cell[     449] = 32'hf6e559db;
    ram_cell[     450] = 32'habec9880;
    ram_cell[     451] = 32'hbad7e88a;
    ram_cell[     452] = 32'hac30e471;
    ram_cell[     453] = 32'h61011f41;
    ram_cell[     454] = 32'h30db5302;
    ram_cell[     455] = 32'h98496e24;
    ram_cell[     456] = 32'h405630b6;
    ram_cell[     457] = 32'ha3cebdec;
    ram_cell[     458] = 32'h58784dcf;
    ram_cell[     459] = 32'hccf95f41;
    ram_cell[     460] = 32'h47e97d15;
    ram_cell[     461] = 32'h624226b2;
    ram_cell[     462] = 32'h2bc01bfb;
    ram_cell[     463] = 32'h5e212b01;
    ram_cell[     464] = 32'hb87b0217;
    ram_cell[     465] = 32'h59a0737c;
    ram_cell[     466] = 32'h7d4a496f;
    ram_cell[     467] = 32'h7ccd4d78;
    ram_cell[     468] = 32'hab027feb;
    ram_cell[     469] = 32'hee91bdff;
    ram_cell[     470] = 32'h9884169f;
    ram_cell[     471] = 32'hea590193;
    ram_cell[     472] = 32'h1e907b25;
    ram_cell[     473] = 32'hdd3b4a0b;
    ram_cell[     474] = 32'h34ed12ed;
    ram_cell[     475] = 32'hefb4ee20;
    ram_cell[     476] = 32'he1b3056c;
    ram_cell[     477] = 32'ha169ee63;
    ram_cell[     478] = 32'h51f6b8d6;
    ram_cell[     479] = 32'h697093e2;
    ram_cell[     480] = 32'h1bbbaf41;
    ram_cell[     481] = 32'hcac2771c;
    ram_cell[     482] = 32'hab6a3455;
    ram_cell[     483] = 32'ha07c5e2c;
    ram_cell[     484] = 32'hc4db6f9d;
    ram_cell[     485] = 32'hc394b652;
    ram_cell[     486] = 32'hd3b1c368;
    ram_cell[     487] = 32'h6f61e417;
    ram_cell[     488] = 32'h5f6db660;
    ram_cell[     489] = 32'h5179fe81;
    ram_cell[     490] = 32'hd164e629;
    ram_cell[     491] = 32'hdbcea628;
    ram_cell[     492] = 32'h58f73f53;
    ram_cell[     493] = 32'hea01b555;
    ram_cell[     494] = 32'h938ac1bc;
    ram_cell[     495] = 32'h83c58054;
    ram_cell[     496] = 32'ha14fcd9e;
    ram_cell[     497] = 32'h86f5f09a;
    ram_cell[     498] = 32'hec842677;
    ram_cell[     499] = 32'h45f2e550;
    ram_cell[     500] = 32'h172b9b57;
    ram_cell[     501] = 32'h8fc9da25;
    ram_cell[     502] = 32'h919b8e28;
    ram_cell[     503] = 32'h796ee5cb;
    ram_cell[     504] = 32'h50c76ddb;
    ram_cell[     505] = 32'hefbfd106;
    ram_cell[     506] = 32'ha94113fc;
    ram_cell[     507] = 32'hf7412c10;
    ram_cell[     508] = 32'h64a43996;
    ram_cell[     509] = 32'ha902a4d3;
    ram_cell[     510] = 32'h0501ad0f;
    ram_cell[     511] = 32'h9e9485e5;
    // src matrix B
    ram_cell[     512] = 32'he3cd1404;
    ram_cell[     513] = 32'h6d74baf3;
    ram_cell[     514] = 32'h1352597b;
    ram_cell[     515] = 32'h770a68c4;
    ram_cell[     516] = 32'hb04d50da;
    ram_cell[     517] = 32'h4bf7b660;
    ram_cell[     518] = 32'h726a0a39;
    ram_cell[     519] = 32'h88fe5110;
    ram_cell[     520] = 32'h863ff721;
    ram_cell[     521] = 32'h73a349d6;
    ram_cell[     522] = 32'h72fdd868;
    ram_cell[     523] = 32'he08ece4e;
    ram_cell[     524] = 32'h9284bd07;
    ram_cell[     525] = 32'h36eb38e6;
    ram_cell[     526] = 32'h3e1b8158;
    ram_cell[     527] = 32'he288414f;
    ram_cell[     528] = 32'hcbb873c5;
    ram_cell[     529] = 32'h2fa79514;
    ram_cell[     530] = 32'h7743c1f7;
    ram_cell[     531] = 32'hfd8e4756;
    ram_cell[     532] = 32'h6e829df1;
    ram_cell[     533] = 32'h64e438ca;
    ram_cell[     534] = 32'h5bb2ddea;
    ram_cell[     535] = 32'h25f0659b;
    ram_cell[     536] = 32'he11a5d85;
    ram_cell[     537] = 32'h499e3d2e;
    ram_cell[     538] = 32'hcebefba7;
    ram_cell[     539] = 32'hb6f2c793;
    ram_cell[     540] = 32'h79a3df4d;
    ram_cell[     541] = 32'h7e7682bd;
    ram_cell[     542] = 32'hde04313d;
    ram_cell[     543] = 32'h45ea55c4;
    ram_cell[     544] = 32'h632d13d6;
    ram_cell[     545] = 32'h86ad9f90;
    ram_cell[     546] = 32'h920e28df;
    ram_cell[     547] = 32'h0405a330;
    ram_cell[     548] = 32'h92a5c5f5;
    ram_cell[     549] = 32'h20ee8c6b;
    ram_cell[     550] = 32'h921668fb;
    ram_cell[     551] = 32'hc5f78f0f;
    ram_cell[     552] = 32'h512ee23b;
    ram_cell[     553] = 32'h544dc3f8;
    ram_cell[     554] = 32'hb6ab54ad;
    ram_cell[     555] = 32'h9bab7c1a;
    ram_cell[     556] = 32'h3d32f58c;
    ram_cell[     557] = 32'hd23be2f0;
    ram_cell[     558] = 32'h52daf96c;
    ram_cell[     559] = 32'h8cdce2ab;
    ram_cell[     560] = 32'h6255f3c9;
    ram_cell[     561] = 32'h5173fc68;
    ram_cell[     562] = 32'h9b24fa81;
    ram_cell[     563] = 32'h58ccfde8;
    ram_cell[     564] = 32'h4a43b13e;
    ram_cell[     565] = 32'he9fc67bc;
    ram_cell[     566] = 32'hc827358b;
    ram_cell[     567] = 32'hacf97e99;
    ram_cell[     568] = 32'h36a63b91;
    ram_cell[     569] = 32'h72faf273;
    ram_cell[     570] = 32'h8d0c6a8d;
    ram_cell[     571] = 32'hf8e21af7;
    ram_cell[     572] = 32'h2090700b;
    ram_cell[     573] = 32'hf75b0bc0;
    ram_cell[     574] = 32'h265f2352;
    ram_cell[     575] = 32'h979a7162;
    ram_cell[     576] = 32'h9c77fccf;
    ram_cell[     577] = 32'he28418a3;
    ram_cell[     578] = 32'h5690abf1;
    ram_cell[     579] = 32'h98f32c53;
    ram_cell[     580] = 32'h42d93be9;
    ram_cell[     581] = 32'h36e8c1bd;
    ram_cell[     582] = 32'h8823eb2c;
    ram_cell[     583] = 32'h4cb1b7e1;
    ram_cell[     584] = 32'h4e26bb67;
    ram_cell[     585] = 32'h40dd4c23;
    ram_cell[     586] = 32'h5237f014;
    ram_cell[     587] = 32'h5015b6cf;
    ram_cell[     588] = 32'hf7781d5d;
    ram_cell[     589] = 32'hb52f5b7d;
    ram_cell[     590] = 32'hf6db65cc;
    ram_cell[     591] = 32'ha6305bda;
    ram_cell[     592] = 32'h5b0f9bee;
    ram_cell[     593] = 32'haef33a80;
    ram_cell[     594] = 32'h0e53c462;
    ram_cell[     595] = 32'hbeadd8c9;
    ram_cell[     596] = 32'h7584c881;
    ram_cell[     597] = 32'h5a044da7;
    ram_cell[     598] = 32'h1811b421;
    ram_cell[     599] = 32'h604f63f4;
    ram_cell[     600] = 32'hbff97503;
    ram_cell[     601] = 32'hc1e333e9;
    ram_cell[     602] = 32'ha0139c17;
    ram_cell[     603] = 32'hbf0175a1;
    ram_cell[     604] = 32'h40d885ce;
    ram_cell[     605] = 32'hec89feae;
    ram_cell[     606] = 32'hfba8287b;
    ram_cell[     607] = 32'hcf090af8;
    ram_cell[     608] = 32'h0c91c306;
    ram_cell[     609] = 32'hcc3120a7;
    ram_cell[     610] = 32'h434dbbc2;
    ram_cell[     611] = 32'h5edab8eb;
    ram_cell[     612] = 32'he66ce99d;
    ram_cell[     613] = 32'h7aeaef65;
    ram_cell[     614] = 32'h6264c33a;
    ram_cell[     615] = 32'hd6369178;
    ram_cell[     616] = 32'h4c8a29f7;
    ram_cell[     617] = 32'he113a8a6;
    ram_cell[     618] = 32'hbde9aed4;
    ram_cell[     619] = 32'hba140888;
    ram_cell[     620] = 32'ha3759fce;
    ram_cell[     621] = 32'hd9d7ae49;
    ram_cell[     622] = 32'he7e72d3f;
    ram_cell[     623] = 32'h24a0a422;
    ram_cell[     624] = 32'hed698dd2;
    ram_cell[     625] = 32'hc289c499;
    ram_cell[     626] = 32'h780a8179;
    ram_cell[     627] = 32'habbbf29b;
    ram_cell[     628] = 32'hc4344b12;
    ram_cell[     629] = 32'h7354e1db;
    ram_cell[     630] = 32'h7c0d81d1;
    ram_cell[     631] = 32'h83527450;
    ram_cell[     632] = 32'h6bded29d;
    ram_cell[     633] = 32'h91853d88;
    ram_cell[     634] = 32'h7cf6eba1;
    ram_cell[     635] = 32'hd57ab043;
    ram_cell[     636] = 32'hcb489b44;
    ram_cell[     637] = 32'hf178a42b;
    ram_cell[     638] = 32'hbd2cf1ee;
    ram_cell[     639] = 32'h23a62381;
    ram_cell[     640] = 32'h5f013836;
    ram_cell[     641] = 32'he29be8f3;
    ram_cell[     642] = 32'h59709ba9;
    ram_cell[     643] = 32'h598d9967;
    ram_cell[     644] = 32'hd2320615;
    ram_cell[     645] = 32'h1add8ebb;
    ram_cell[     646] = 32'hab9beda2;
    ram_cell[     647] = 32'h47a0995b;
    ram_cell[     648] = 32'h717bab85;
    ram_cell[     649] = 32'hab7439ac;
    ram_cell[     650] = 32'h632832a5;
    ram_cell[     651] = 32'h44473790;
    ram_cell[     652] = 32'h713f6f00;
    ram_cell[     653] = 32'h2a5c42ef;
    ram_cell[     654] = 32'he8365b49;
    ram_cell[     655] = 32'hc60ecd08;
    ram_cell[     656] = 32'h836891bf;
    ram_cell[     657] = 32'h4cff689a;
    ram_cell[     658] = 32'h9964b69e;
    ram_cell[     659] = 32'h4e3ebb65;
    ram_cell[     660] = 32'hd46029ca;
    ram_cell[     661] = 32'h242bcf57;
    ram_cell[     662] = 32'he5e8ee02;
    ram_cell[     663] = 32'h1dc45237;
    ram_cell[     664] = 32'hdea6abf9;
    ram_cell[     665] = 32'h53493bf7;
    ram_cell[     666] = 32'h1764d9c1;
    ram_cell[     667] = 32'hbaeb537c;
    ram_cell[     668] = 32'hace0e173;
    ram_cell[     669] = 32'h02c98715;
    ram_cell[     670] = 32'h6c1ea80f;
    ram_cell[     671] = 32'hd86c2660;
    ram_cell[     672] = 32'h7c07eea2;
    ram_cell[     673] = 32'h20440233;
    ram_cell[     674] = 32'h7914ca91;
    ram_cell[     675] = 32'hf2ed7c2b;
    ram_cell[     676] = 32'h0a10e0c6;
    ram_cell[     677] = 32'h552a12c8;
    ram_cell[     678] = 32'h4ad947ec;
    ram_cell[     679] = 32'he289f2b7;
    ram_cell[     680] = 32'h9952189f;
    ram_cell[     681] = 32'hd59aca46;
    ram_cell[     682] = 32'h4216fae1;
    ram_cell[     683] = 32'h0cae2ac2;
    ram_cell[     684] = 32'h75862cde;
    ram_cell[     685] = 32'hceaedd83;
    ram_cell[     686] = 32'hb692aabd;
    ram_cell[     687] = 32'hbe52a381;
    ram_cell[     688] = 32'h6ffb0d42;
    ram_cell[     689] = 32'h654e8cbb;
    ram_cell[     690] = 32'h9309273d;
    ram_cell[     691] = 32'h66ba1458;
    ram_cell[     692] = 32'hc0c2f150;
    ram_cell[     693] = 32'hb7c77845;
    ram_cell[     694] = 32'h0374232c;
    ram_cell[     695] = 32'ha72a250a;
    ram_cell[     696] = 32'hc51081d1;
    ram_cell[     697] = 32'h374b6ecb;
    ram_cell[     698] = 32'h2ff6f54d;
    ram_cell[     699] = 32'h6a9252c4;
    ram_cell[     700] = 32'hcf35001c;
    ram_cell[     701] = 32'h1688903e;
    ram_cell[     702] = 32'h975aa69a;
    ram_cell[     703] = 32'h6b675d17;
    ram_cell[     704] = 32'hdab456da;
    ram_cell[     705] = 32'he582061e;
    ram_cell[     706] = 32'h61996ec7;
    ram_cell[     707] = 32'h22ffe374;
    ram_cell[     708] = 32'h77f281bb;
    ram_cell[     709] = 32'h0acf1620;
    ram_cell[     710] = 32'h754ec90d;
    ram_cell[     711] = 32'ha2ccf948;
    ram_cell[     712] = 32'h1a40c069;
    ram_cell[     713] = 32'hded3b080;
    ram_cell[     714] = 32'h2068f136;
    ram_cell[     715] = 32'he87b21c7;
    ram_cell[     716] = 32'hf9ef834b;
    ram_cell[     717] = 32'h498ddbb3;
    ram_cell[     718] = 32'hbd2991ea;
    ram_cell[     719] = 32'h3d23d5dc;
    ram_cell[     720] = 32'ha738dbe3;
    ram_cell[     721] = 32'h01480993;
    ram_cell[     722] = 32'h862bc745;
    ram_cell[     723] = 32'h27764144;
    ram_cell[     724] = 32'h90fa0579;
    ram_cell[     725] = 32'hc8093ff8;
    ram_cell[     726] = 32'hac9b9fdd;
    ram_cell[     727] = 32'h2a786e64;
    ram_cell[     728] = 32'ha062a735;
    ram_cell[     729] = 32'hbfa9f88e;
    ram_cell[     730] = 32'h46258620;
    ram_cell[     731] = 32'h06bd104a;
    ram_cell[     732] = 32'h7e85cb72;
    ram_cell[     733] = 32'h3886e200;
    ram_cell[     734] = 32'h4962d144;
    ram_cell[     735] = 32'hc1be98bc;
    ram_cell[     736] = 32'h11b26ba0;
    ram_cell[     737] = 32'h7abd4b60;
    ram_cell[     738] = 32'h59ca2904;
    ram_cell[     739] = 32'h148cfa94;
    ram_cell[     740] = 32'h4acaf6e4;
    ram_cell[     741] = 32'hb5888132;
    ram_cell[     742] = 32'h6cef3d44;
    ram_cell[     743] = 32'h9b6a466f;
    ram_cell[     744] = 32'hab4b9438;
    ram_cell[     745] = 32'hc6affe34;
    ram_cell[     746] = 32'h580e15ef;
    ram_cell[     747] = 32'hb5a81262;
    ram_cell[     748] = 32'hc61f19b5;
    ram_cell[     749] = 32'h058ead96;
    ram_cell[     750] = 32'he929b051;
    ram_cell[     751] = 32'h25d0b363;
    ram_cell[     752] = 32'hc2479cdd;
    ram_cell[     753] = 32'ha3d0b660;
    ram_cell[     754] = 32'hbcf9f9ee;
    ram_cell[     755] = 32'hf151c987;
    ram_cell[     756] = 32'h3a768fac;
    ram_cell[     757] = 32'h6fd43d98;
    ram_cell[     758] = 32'h2282204d;
    ram_cell[     759] = 32'h40d4e870;
    ram_cell[     760] = 32'h173f6a8c;
    ram_cell[     761] = 32'h840d29e7;
    ram_cell[     762] = 32'h64298050;
    ram_cell[     763] = 32'hb7343564;
    ram_cell[     764] = 32'h12a460d6;
    ram_cell[     765] = 32'hcad3a29b;
    ram_cell[     766] = 32'hb5b9a863;
    ram_cell[     767] = 32'h52fc5dc8;
end

endmodule

