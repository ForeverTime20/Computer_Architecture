
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

//qsort
// initial begin
//     // qsort 256
//     ram_cell[       0] = 32'h0000009a;
//     ram_cell[       1] = 32'h000000e3;
//     ram_cell[       2] = 32'h0000002b;
//     ram_cell[       3] = 32'h0000001c;
//     ram_cell[       4] = 32'h00000074;
//     ram_cell[       5] = 32'h00000091;
//     ram_cell[       6] = 32'h0000007b;
//     ram_cell[       7] = 32'h000000aa;
//     ram_cell[       8] = 32'h00000073;
//     ram_cell[       9] = 32'h000000ae;
//     ram_cell[      10] = 32'h00000069;
//     ram_cell[      11] = 32'h00000097;
//     ram_cell[      12] = 32'h00000098;
//     ram_cell[      13] = 32'h000000c1;
//     ram_cell[      14] = 32'h00000030;
//     ram_cell[      15] = 32'h00000047;
//     ram_cell[      16] = 32'h0000002c;
//     ram_cell[      17] = 32'h000000d8;
//     ram_cell[      18] = 32'h000000f8;
//     ram_cell[      19] = 32'h00000034;
//     ram_cell[      20] = 32'h0000005d;
//     ram_cell[      21] = 32'h0000006e;
//     ram_cell[      22] = 32'h0000007f;
//     ram_cell[      23] = 32'h000000a8;
//     ram_cell[      24] = 32'h000000b0;
//     ram_cell[      25] = 32'h000000e0;
//     ram_cell[      26] = 32'h000000f2;
//     ram_cell[      27] = 32'h00000095;
//     ram_cell[      28] = 32'h00000066;
//     ram_cell[      29] = 32'h00000053;
//     ram_cell[      30] = 32'h00000035;
//     ram_cell[      31] = 32'h000000da;
//     ram_cell[      32] = 32'h00000094;
//     ram_cell[      33] = 32'h000000b7;
//     ram_cell[      34] = 32'h00000019;
//     ram_cell[      35] = 32'h000000d1;
//     ram_cell[      36] = 32'h0000008e;
//     ram_cell[      37] = 32'h00000057;
//     ram_cell[      38] = 32'h0000003a;
//     ram_cell[      39] = 32'h000000c7;
//     ram_cell[      40] = 32'h0000006f;
//     ram_cell[      41] = 32'h000000d3;
//     ram_cell[      42] = 32'h000000d4;
//     ram_cell[      43] = 32'h00000085;
//     ram_cell[      44] = 32'h000000cd;
//     ram_cell[      45] = 32'h000000dc;
//     ram_cell[      46] = 32'h00000003;
//     ram_cell[      47] = 32'h0000009f;
//     ram_cell[      48] = 32'h0000007c;
//     ram_cell[      49] = 32'h0000005a;
//     ram_cell[      50] = 32'h00000093;
//     ram_cell[      51] = 32'h000000de;
//     ram_cell[      52] = 32'h0000000c;
//     ram_cell[      53] = 32'h000000d2;
//     ram_cell[      54] = 32'h0000006d;
//     ram_cell[      55] = 32'h0000002e;
//     ram_cell[      56] = 32'h000000df;
//     ram_cell[      57] = 32'h0000003c;
//     ram_cell[      58] = 32'h00000072;
//     ram_cell[      59] = 32'h000000f4;
//     ram_cell[      60] = 32'h0000004c;
//     ram_cell[      61] = 32'h00000079;
//     ram_cell[      62] = 32'h00000016;
//     ram_cell[      63] = 32'h00000028;
//     ram_cell[      64] = 32'h00000054;
//     ram_cell[      65] = 32'h0000003d;
//     ram_cell[      66] = 32'h000000ba;
//     ram_cell[      67] = 32'h000000b1;
//     ram_cell[      68] = 32'h000000c3;
//     ram_cell[      69] = 32'h0000008a;
//     ram_cell[      70] = 32'h0000008c;
//     ram_cell[      71] = 32'h000000cb;
//     ram_cell[      72] = 32'h00000081;
//     ram_cell[      73] = 32'h0000009c;
//     ram_cell[      74] = 32'h0000002f;
//     ram_cell[      75] = 32'h000000b2;
//     ram_cell[      76] = 32'h00000027;
//     ram_cell[      77] = 32'h00000031;
//     ram_cell[      78] = 32'h00000082;
//     ram_cell[      79] = 32'h00000086;
//     ram_cell[      80] = 32'h00000092;
//     ram_cell[      81] = 32'h000000e1;
//     ram_cell[      82] = 32'h00000037;
//     ram_cell[      83] = 32'h00000075;
//     ram_cell[      84] = 32'h0000000f;
//     ram_cell[      85] = 32'h000000c2;
//     ram_cell[      86] = 32'h00000044;
//     ram_cell[      87] = 32'h0000004d;
//     ram_cell[      88] = 32'h00000062;
//     ram_cell[      89] = 32'h000000b4;
//     ram_cell[      90] = 32'h000000af;
//     ram_cell[      91] = 32'h0000001e;
//     ram_cell[      92] = 32'h00000012;
//     ram_cell[      93] = 32'h000000a9;
//     ram_cell[      94] = 32'h000000d0;
//     ram_cell[      95] = 32'h000000b9;
//     ram_cell[      96] = 32'h0000007d;
//     ram_cell[      97] = 32'h00000040;
//     ram_cell[      98] = 32'h00000007;
//     ram_cell[      99] = 32'h000000a2;
//     ram_cell[     100] = 32'h000000ca;
//     ram_cell[     101] = 32'h0000006b;
//     ram_cell[     102] = 32'h00000052;
//     ram_cell[     103] = 32'h000000c5;
//     ram_cell[     104] = 32'h000000d9;
//     ram_cell[     105] = 32'h00000002;
//     ram_cell[     106] = 32'h000000ac;
//     ram_cell[     107] = 32'h0000000b;
//     ram_cell[     108] = 32'h0000007e;
//     ram_cell[     109] = 32'h00000061;
//     ram_cell[     110] = 32'h00000068;
//     ram_cell[     111] = 32'h000000fb;
//     ram_cell[     112] = 32'h0000004a;
//     ram_cell[     113] = 32'h000000a0;
//     ram_cell[     114] = 32'h000000e7;
//     ram_cell[     115] = 32'h00000049;
//     ram_cell[     116] = 32'h00000013;
//     ram_cell[     117] = 32'h00000032;
//     ram_cell[     118] = 32'h000000b5;
//     ram_cell[     119] = 32'h00000080;
//     ram_cell[     120] = 32'h00000077;
//     ram_cell[     121] = 32'h00000001;
//     ram_cell[     122] = 32'h0000008f;
//     ram_cell[     123] = 32'h0000000d;
//     ram_cell[     124] = 32'h0000009e;
//     ram_cell[     125] = 32'h000000ea;
//     ram_cell[     126] = 32'h0000001b;
//     ram_cell[     127] = 32'h000000b6;
//     ram_cell[     128] = 32'h0000006a;
//     ram_cell[     129] = 32'h000000e5;
//     ram_cell[     130] = 32'h00000014;
//     ram_cell[     131] = 32'h000000e8;
//     ram_cell[     132] = 32'h00000078;
//     ram_cell[     133] = 32'h00000084;
//     ram_cell[     134] = 32'h000000ef;
//     ram_cell[     135] = 32'h00000046;
//     ram_cell[     136] = 32'h000000f9;
//     ram_cell[     137] = 32'h00000063;
//     ram_cell[     138] = 32'h0000001d;
//     ram_cell[     139] = 32'h0000005c;
//     ram_cell[     140] = 32'h00000018;
//     ram_cell[     141] = 32'h000000bc;
//     ram_cell[     142] = 32'h000000ee;
//     ram_cell[     143] = 32'h00000005;
//     ram_cell[     144] = 32'h00000045;
//     ram_cell[     145] = 32'h00000021;
//     ram_cell[     146] = 32'h000000e6;
//     ram_cell[     147] = 32'h000000ed;
//     ram_cell[     148] = 32'h000000fa;
//     ram_cell[     149] = 32'h000000db;
//     ram_cell[     150] = 32'h00000011;
//     ram_cell[     151] = 32'h00000065;
//     ram_cell[     152] = 32'h00000009;
//     ram_cell[     153] = 32'h000000b8;
//     ram_cell[     154] = 32'h00000024;
//     ram_cell[     155] = 32'h00000096;
//     ram_cell[     156] = 32'h00000071;
//     ram_cell[     157] = 32'h00000048;
//     ram_cell[     158] = 32'h0000003e;
//     ram_cell[     159] = 32'h0000007a;
//     ram_cell[     160] = 32'h000000f5;
//     ram_cell[     161] = 32'h00000067;
//     ram_cell[     162] = 32'h000000bf;
//     ram_cell[     163] = 32'h000000f1;
//     ram_cell[     164] = 32'h00000055;
//     ram_cell[     165] = 32'h000000ff;
//     ram_cell[     166] = 32'h00000042;
//     ram_cell[     167] = 32'h000000b3;
//     ram_cell[     168] = 32'h00000020;
//     ram_cell[     169] = 32'h000000fd;
//     ram_cell[     170] = 32'h000000a6;
//     ram_cell[     171] = 32'h00000064;
//     ram_cell[     172] = 32'h0000005f;
//     ram_cell[     173] = 32'h000000ab;
//     ram_cell[     174] = 32'h000000fe;
//     ram_cell[     175] = 32'h000000c9;
//     ram_cell[     176] = 32'h000000dd;
//     ram_cell[     177] = 32'h00000043;
//     ram_cell[     178] = 32'h00000025;
//     ram_cell[     179] = 32'h000000a5;
//     ram_cell[     180] = 32'h0000000a;
//     ram_cell[     181] = 32'h0000005b;
//     ram_cell[     182] = 32'h0000001a;
//     ram_cell[     183] = 32'h000000bb;
//     ram_cell[     184] = 32'h0000006c;
//     ram_cell[     185] = 32'h000000cc;
//     ram_cell[     186] = 32'h00000023;
//     ram_cell[     187] = 32'h00000076;
//     ram_cell[     188] = 32'h0000004f;
//     ram_cell[     189] = 32'h000000be;
//     ram_cell[     190] = 32'h00000029;
//     ram_cell[     191] = 32'h00000083;
//     ram_cell[     192] = 32'h0000002a;
//     ram_cell[     193] = 32'h000000fc;
//     ram_cell[     194] = 32'h00000026;
//     ram_cell[     195] = 32'h00000038;
//     ram_cell[     196] = 32'h0000000e;
//     ram_cell[     197] = 32'h000000ce;
//     ram_cell[     198] = 32'h00000036;
//     ram_cell[     199] = 32'h00000015;
//     ram_cell[     200] = 32'h00000056;
//     ram_cell[     201] = 32'h0000009b;
//     ram_cell[     202] = 32'h00000059;
//     ram_cell[     203] = 32'h00000090;
//     ram_cell[     204] = 32'h000000d5;
//     ram_cell[     205] = 32'h0000009d;
//     ram_cell[     206] = 32'h000000c4;
//     ram_cell[     207] = 32'h000000ad;
//     ram_cell[     208] = 32'h0000002d;
//     ram_cell[     209] = 32'h000000a7;
//     ram_cell[     210] = 32'h000000cf;
//     ram_cell[     211] = 32'h00000010;
//     ram_cell[     212] = 32'h00000058;
//     ram_cell[     213] = 32'h00000022;
//     ram_cell[     214] = 32'h00000000;
//     ram_cell[     215] = 32'h000000d7;
//     ram_cell[     216] = 32'h00000039;
//     ram_cell[     217] = 32'h00000008;
//     ram_cell[     218] = 32'h000000c0;
//     ram_cell[     219] = 32'h00000087;
//     ram_cell[     220] = 32'h000000bd;
//     ram_cell[     221] = 32'h00000006;
//     ram_cell[     222] = 32'h0000005e;
//     ram_cell[     223] = 32'h000000eb;
//     ram_cell[     224] = 32'h000000ec;
//     ram_cell[     225] = 32'h00000060;
//     ram_cell[     226] = 32'h000000a3;
//     ram_cell[     227] = 32'h000000c8;
//     ram_cell[     228] = 32'h00000089;
//     ram_cell[     229] = 32'h0000004b;
//     ram_cell[     230] = 32'h000000c6;
//     ram_cell[     231] = 32'h0000003b;
//     ram_cell[     232] = 32'h000000a4;
//     ram_cell[     233] = 32'h000000f3;
//     ram_cell[     234] = 32'h00000004;
//     ram_cell[     235] = 32'h000000f6;
//     ram_cell[     236] = 32'h000000a1;
//     ram_cell[     237] = 32'h00000070;
//     ram_cell[     238] = 32'h000000f0;
//     ram_cell[     239] = 32'h000000e4;
//     ram_cell[     240] = 32'h000000f7;
//     ram_cell[     241] = 32'h00000033;
//     ram_cell[     242] = 32'h0000008b;
//     ram_cell[     243] = 32'h000000e9;
//     ram_cell[     244] = 32'h0000003f;
//     ram_cell[     245] = 32'h0000008d;
//     ram_cell[     246] = 32'h000000e2;
//     ram_cell[     247] = 32'h00000041;
//     ram_cell[     248] = 32'h00000017;
//     ram_cell[     249] = 32'h0000004e;
//     ram_cell[     250] = 32'h0000001f;
//     ram_cell[     251] = 32'h00000088;
//     ram_cell[     252] = 32'h000000d6;
//     ram_cell[     253] = 32'h00000050;
//     ram_cell[     254] = 32'h00000099;
//     ram_cell[     255] = 32'h00000051;
// end

//matrix
initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'h791fcd2e;
    ram_cell[       1] = 32'h0;  // 32'heff3d520;
    ram_cell[       2] = 32'h0;  // 32'hbd847b84;
    ram_cell[       3] = 32'h0;  // 32'hb0e9c84b;
    ram_cell[       4] = 32'h0;  // 32'h38570320;
    ram_cell[       5] = 32'h0;  // 32'hbb76e841;
    ram_cell[       6] = 32'h0;  // 32'h224f2629;
    ram_cell[       7] = 32'h0;  // 32'h1ebf2170;
    ram_cell[       8] = 32'h0;  // 32'hd7b5f3db;
    ram_cell[       9] = 32'h0;  // 32'h5ee57156;
    ram_cell[      10] = 32'h0;  // 32'hf9c8be7f;
    ram_cell[      11] = 32'h0;  // 32'h4ba07f20;
    ram_cell[      12] = 32'h0;  // 32'h1d67393d;
    ram_cell[      13] = 32'h0;  // 32'h48d7e735;
    ram_cell[      14] = 32'h0;  // 32'h62aaf7b7;
    ram_cell[      15] = 32'h0;  // 32'hd8673717;
    ram_cell[      16] = 32'h0;  // 32'hc9c91a84;
    ram_cell[      17] = 32'h0;  // 32'h8ba26243;
    ram_cell[      18] = 32'h0;  // 32'h1959f638;
    ram_cell[      19] = 32'h0;  // 32'hdb632495;
    ram_cell[      20] = 32'h0;  // 32'h59ebccd5;
    ram_cell[      21] = 32'h0;  // 32'h202af67b;
    ram_cell[      22] = 32'h0;  // 32'h5f52f300;
    ram_cell[      23] = 32'h0;  // 32'h00ce2b2a;
    ram_cell[      24] = 32'h0;  // 32'h9d501e8d;
    ram_cell[      25] = 32'h0;  // 32'h5c36d6e9;
    ram_cell[      26] = 32'h0;  // 32'h765e7502;
    ram_cell[      27] = 32'h0;  // 32'h50b8a7bd;
    ram_cell[      28] = 32'h0;  // 32'hbc540ad7;
    ram_cell[      29] = 32'h0;  // 32'h8894899d;
    ram_cell[      30] = 32'h0;  // 32'hfb067457;
    ram_cell[      31] = 32'h0;  // 32'hdf17e924;
    ram_cell[      32] = 32'h0;  // 32'h219b411f;
    ram_cell[      33] = 32'h0;  // 32'hcfdd38fa;
    ram_cell[      34] = 32'h0;  // 32'hcde05e82;
    ram_cell[      35] = 32'h0;  // 32'h54b16638;
    ram_cell[      36] = 32'h0;  // 32'h9447d112;
    ram_cell[      37] = 32'h0;  // 32'hb4760b24;
    ram_cell[      38] = 32'h0;  // 32'ha9fcf8be;
    ram_cell[      39] = 32'h0;  // 32'h3b434282;
    ram_cell[      40] = 32'h0;  // 32'h108fc785;
    ram_cell[      41] = 32'h0;  // 32'hd1d5cced;
    ram_cell[      42] = 32'h0;  // 32'h7041655d;
    ram_cell[      43] = 32'h0;  // 32'hf5ab90d0;
    ram_cell[      44] = 32'h0;  // 32'h57b61cda;
    ram_cell[      45] = 32'h0;  // 32'h13195141;
    ram_cell[      46] = 32'h0;  // 32'h735ba45f;
    ram_cell[      47] = 32'h0;  // 32'haf8c542c;
    ram_cell[      48] = 32'h0;  // 32'hc9d6981a;
    ram_cell[      49] = 32'h0;  // 32'h03a33c11;
    ram_cell[      50] = 32'h0;  // 32'h1b003227;
    ram_cell[      51] = 32'h0;  // 32'hc278d121;
    ram_cell[      52] = 32'h0;  // 32'h4e7ce87d;
    ram_cell[      53] = 32'h0;  // 32'hf4bc2fd2;
    ram_cell[      54] = 32'h0;  // 32'h68e180f3;
    ram_cell[      55] = 32'h0;  // 32'h0d5c9151;
    ram_cell[      56] = 32'h0;  // 32'ha0ef55cf;
    ram_cell[      57] = 32'h0;  // 32'hf28e8db9;
    ram_cell[      58] = 32'h0;  // 32'h0f55e23f;
    ram_cell[      59] = 32'h0;  // 32'h17e39cc4;
    ram_cell[      60] = 32'h0;  // 32'h1ccf145c;
    ram_cell[      61] = 32'h0;  // 32'hded473b6;
    ram_cell[      62] = 32'h0;  // 32'h4b9ce2f9;
    ram_cell[      63] = 32'h0;  // 32'hfc8a4e3e;
    ram_cell[      64] = 32'h0;  // 32'h1ee60a4b;
    ram_cell[      65] = 32'h0;  // 32'hd7f35d8d;
    ram_cell[      66] = 32'h0;  // 32'h8b1157e7;
    ram_cell[      67] = 32'h0;  // 32'h89eb2466;
    ram_cell[      68] = 32'h0;  // 32'hfee7c73f;
    ram_cell[      69] = 32'h0;  // 32'hf4c4e993;
    ram_cell[      70] = 32'h0;  // 32'h544cb15f;
    ram_cell[      71] = 32'h0;  // 32'h33d31990;
    ram_cell[      72] = 32'h0;  // 32'h7ffbddab;
    ram_cell[      73] = 32'h0;  // 32'h1245e393;
    ram_cell[      74] = 32'h0;  // 32'h090d5eb7;
    ram_cell[      75] = 32'h0;  // 32'haa951c62;
    ram_cell[      76] = 32'h0;  // 32'h09f13df5;
    ram_cell[      77] = 32'h0;  // 32'hdbc3b50a;
    ram_cell[      78] = 32'h0;  // 32'hc28adf76;
    ram_cell[      79] = 32'h0;  // 32'hcb437a61;
    ram_cell[      80] = 32'h0;  // 32'h09538767;
    ram_cell[      81] = 32'h0;  // 32'h5b807965;
    ram_cell[      82] = 32'h0;  // 32'hf79966ee;
    ram_cell[      83] = 32'h0;  // 32'ha39a1897;
    ram_cell[      84] = 32'h0;  // 32'h5fae9922;
    ram_cell[      85] = 32'h0;  // 32'h7e28acdb;
    ram_cell[      86] = 32'h0;  // 32'h5cd5043d;
    ram_cell[      87] = 32'h0;  // 32'h7b904fe5;
    ram_cell[      88] = 32'h0;  // 32'h7e02c10d;
    ram_cell[      89] = 32'h0;  // 32'h0506b879;
    ram_cell[      90] = 32'h0;  // 32'he2c90585;
    ram_cell[      91] = 32'h0;  // 32'h43c7a1fd;
    ram_cell[      92] = 32'h0;  // 32'hdb09895a;
    ram_cell[      93] = 32'h0;  // 32'h81ac519b;
    ram_cell[      94] = 32'h0;  // 32'h851ed5d1;
    ram_cell[      95] = 32'h0;  // 32'h486813e5;
    ram_cell[      96] = 32'h0;  // 32'hafb8aa71;
    ram_cell[      97] = 32'h0;  // 32'h2f5c69c9;
    ram_cell[      98] = 32'h0;  // 32'h4809314c;
    ram_cell[      99] = 32'h0;  // 32'h4e7959bb;
    ram_cell[     100] = 32'h0;  // 32'h222d59e4;
    ram_cell[     101] = 32'h0;  // 32'h4feaf83a;
    ram_cell[     102] = 32'h0;  // 32'h1f207800;
    ram_cell[     103] = 32'h0;  // 32'hcf3048c0;
    ram_cell[     104] = 32'h0;  // 32'h89388af6;
    ram_cell[     105] = 32'h0;  // 32'h44415086;
    ram_cell[     106] = 32'h0;  // 32'hcd24f5d5;
    ram_cell[     107] = 32'h0;  // 32'h51cbeaa6;
    ram_cell[     108] = 32'h0;  // 32'he0922539;
    ram_cell[     109] = 32'h0;  // 32'h59d44e7b;
    ram_cell[     110] = 32'h0;  // 32'h555cf4a9;
    ram_cell[     111] = 32'h0;  // 32'h2d6c7675;
    ram_cell[     112] = 32'h0;  // 32'h87cb6312;
    ram_cell[     113] = 32'h0;  // 32'h6d8f4129;
    ram_cell[     114] = 32'h0;  // 32'h580be921;
    ram_cell[     115] = 32'h0;  // 32'hef6b52c4;
    ram_cell[     116] = 32'h0;  // 32'hc0987ca9;
    ram_cell[     117] = 32'h0;  // 32'h12625980;
    ram_cell[     118] = 32'h0;  // 32'h62c1f7c6;
    ram_cell[     119] = 32'h0;  // 32'hf5e2a4d5;
    ram_cell[     120] = 32'h0;  // 32'hec5283ec;
    ram_cell[     121] = 32'h0;  // 32'h846a1108;
    ram_cell[     122] = 32'h0;  // 32'h548ab196;
    ram_cell[     123] = 32'h0;  // 32'h8c2b67ff;
    ram_cell[     124] = 32'h0;  // 32'h4377389f;
    ram_cell[     125] = 32'h0;  // 32'ha488bb0e;
    ram_cell[     126] = 32'h0;  // 32'h0b763cb3;
    ram_cell[     127] = 32'h0;  // 32'h42df7932;
    ram_cell[     128] = 32'h0;  // 32'hfd702511;
    ram_cell[     129] = 32'h0;  // 32'h725e1a4c;
    ram_cell[     130] = 32'h0;  // 32'hc53621f7;
    ram_cell[     131] = 32'h0;  // 32'h481d0db2;
    ram_cell[     132] = 32'h0;  // 32'h4fb97212;
    ram_cell[     133] = 32'h0;  // 32'h892d120b;
    ram_cell[     134] = 32'h0;  // 32'hf0f72695;
    ram_cell[     135] = 32'h0;  // 32'h1a7a7a56;
    ram_cell[     136] = 32'h0;  // 32'h9fe7d3de;
    ram_cell[     137] = 32'h0;  // 32'hf3cceac0;
    ram_cell[     138] = 32'h0;  // 32'h7e7c1159;
    ram_cell[     139] = 32'h0;  // 32'h211ef327;
    ram_cell[     140] = 32'h0;  // 32'he87d30de;
    ram_cell[     141] = 32'h0;  // 32'h1d2c0188;
    ram_cell[     142] = 32'h0;  // 32'he062d453;
    ram_cell[     143] = 32'h0;  // 32'h532cbb0d;
    ram_cell[     144] = 32'h0;  // 32'ha907718f;
    ram_cell[     145] = 32'h0;  // 32'hd0bb92f7;
    ram_cell[     146] = 32'h0;  // 32'h3f8af532;
    ram_cell[     147] = 32'h0;  // 32'hbf222faf;
    ram_cell[     148] = 32'h0;  // 32'h11970723;
    ram_cell[     149] = 32'h0;  // 32'he4f25d9e;
    ram_cell[     150] = 32'h0;  // 32'h830ca25b;
    ram_cell[     151] = 32'h0;  // 32'h31b3dfb7;
    ram_cell[     152] = 32'h0;  // 32'hc5d231cb;
    ram_cell[     153] = 32'h0;  // 32'h072a50b1;
    ram_cell[     154] = 32'h0;  // 32'h8b1708b4;
    ram_cell[     155] = 32'h0;  // 32'h790b813f;
    ram_cell[     156] = 32'h0;  // 32'h81dd2251;
    ram_cell[     157] = 32'h0;  // 32'hc4b42c97;
    ram_cell[     158] = 32'h0;  // 32'hfded9c7f;
    ram_cell[     159] = 32'h0;  // 32'hc61ba6ab;
    ram_cell[     160] = 32'h0;  // 32'hef806fec;
    ram_cell[     161] = 32'h0;  // 32'h6ada293c;
    ram_cell[     162] = 32'h0;  // 32'h9b7d50bd;
    ram_cell[     163] = 32'h0;  // 32'hcd83c24c;
    ram_cell[     164] = 32'h0;  // 32'hca14f2be;
    ram_cell[     165] = 32'h0;  // 32'ha6dfdbae;
    ram_cell[     166] = 32'h0;  // 32'h013b3b48;
    ram_cell[     167] = 32'h0;  // 32'hdd43f8ff;
    ram_cell[     168] = 32'h0;  // 32'h985d99e3;
    ram_cell[     169] = 32'h0;  // 32'h7968de09;
    ram_cell[     170] = 32'h0;  // 32'h08a5455f;
    ram_cell[     171] = 32'h0;  // 32'h605014b7;
    ram_cell[     172] = 32'h0;  // 32'ha3df9e3c;
    ram_cell[     173] = 32'h0;  // 32'h1797a6eb;
    ram_cell[     174] = 32'h0;  // 32'h84afb8d0;
    ram_cell[     175] = 32'h0;  // 32'h2fbccacd;
    ram_cell[     176] = 32'h0;  // 32'h782b9d46;
    ram_cell[     177] = 32'h0;  // 32'hf59cc159;
    ram_cell[     178] = 32'h0;  // 32'h8b4cba86;
    ram_cell[     179] = 32'h0;  // 32'hc86dfa86;
    ram_cell[     180] = 32'h0;  // 32'h3c29e2fe;
    ram_cell[     181] = 32'h0;  // 32'h96b10bb5;
    ram_cell[     182] = 32'h0;  // 32'h0f12b2f0;
    ram_cell[     183] = 32'h0;  // 32'h9c45f5e3;
    ram_cell[     184] = 32'h0;  // 32'hc7bd441b;
    ram_cell[     185] = 32'h0;  // 32'h228df2e4;
    ram_cell[     186] = 32'h0;  // 32'hfe06cc42;
    ram_cell[     187] = 32'h0;  // 32'he6e61944;
    ram_cell[     188] = 32'h0;  // 32'h6c8bf27f;
    ram_cell[     189] = 32'h0;  // 32'h0c3f254c;
    ram_cell[     190] = 32'h0;  // 32'ha3a076c0;
    ram_cell[     191] = 32'h0;  // 32'h94a32867;
    ram_cell[     192] = 32'h0;  // 32'h2c1256cc;
    ram_cell[     193] = 32'h0;  // 32'hf8c23655;
    ram_cell[     194] = 32'h0;  // 32'hc0542716;
    ram_cell[     195] = 32'h0;  // 32'h95a7f5bd;
    ram_cell[     196] = 32'h0;  // 32'h81c37b99;
    ram_cell[     197] = 32'h0;  // 32'h02110573;
    ram_cell[     198] = 32'h0;  // 32'ha2276c4b;
    ram_cell[     199] = 32'h0;  // 32'h83424132;
    ram_cell[     200] = 32'h0;  // 32'hb3bed909;
    ram_cell[     201] = 32'h0;  // 32'he54b83a8;
    ram_cell[     202] = 32'h0;  // 32'hf32bce79;
    ram_cell[     203] = 32'h0;  // 32'h0fe32769;
    ram_cell[     204] = 32'h0;  // 32'hd289cb24;
    ram_cell[     205] = 32'h0;  // 32'hac98d578;
    ram_cell[     206] = 32'h0;  // 32'hd1f661e1;
    ram_cell[     207] = 32'h0;  // 32'hc4fc79d2;
    ram_cell[     208] = 32'h0;  // 32'h2c0bc621;
    ram_cell[     209] = 32'h0;  // 32'h6b777400;
    ram_cell[     210] = 32'h0;  // 32'h8551921e;
    ram_cell[     211] = 32'h0;  // 32'h3c510a8f;
    ram_cell[     212] = 32'h0;  // 32'habe37f18;
    ram_cell[     213] = 32'h0;  // 32'hae439c37;
    ram_cell[     214] = 32'h0;  // 32'h5146fda5;
    ram_cell[     215] = 32'h0;  // 32'hbdeae054;
    ram_cell[     216] = 32'h0;  // 32'h88ad83b7;
    ram_cell[     217] = 32'h0;  // 32'h884eff75;
    ram_cell[     218] = 32'h0;  // 32'h041c1729;
    ram_cell[     219] = 32'h0;  // 32'hd051a747;
    ram_cell[     220] = 32'h0;  // 32'h53298017;
    ram_cell[     221] = 32'h0;  // 32'heaf9a6e0;
    ram_cell[     222] = 32'h0;  // 32'hf85fa621;
    ram_cell[     223] = 32'h0;  // 32'h4b7ba8f5;
    ram_cell[     224] = 32'h0;  // 32'h9d5a1b71;
    ram_cell[     225] = 32'h0;  // 32'h25cd2ddf;
    ram_cell[     226] = 32'h0;  // 32'h7da820af;
    ram_cell[     227] = 32'h0;  // 32'h5d27daee;
    ram_cell[     228] = 32'h0;  // 32'h451b10bd;
    ram_cell[     229] = 32'h0;  // 32'hb5d75725;
    ram_cell[     230] = 32'h0;  // 32'h491eca7f;
    ram_cell[     231] = 32'h0;  // 32'h5880b39c;
    ram_cell[     232] = 32'h0;  // 32'h782fb04d;
    ram_cell[     233] = 32'h0;  // 32'h438cf65f;
    ram_cell[     234] = 32'h0;  // 32'hc1fc7560;
    ram_cell[     235] = 32'h0;  // 32'hd72979f0;
    ram_cell[     236] = 32'h0;  // 32'hc5e0510d;
    ram_cell[     237] = 32'h0;  // 32'he6971bee;
    ram_cell[     238] = 32'h0;  // 32'heb17390f;
    ram_cell[     239] = 32'h0;  // 32'h980adf5b;
    ram_cell[     240] = 32'h0;  // 32'h0acdfb6f;
    ram_cell[     241] = 32'h0;  // 32'h1363808b;
    ram_cell[     242] = 32'h0;  // 32'h417f477d;
    ram_cell[     243] = 32'h0;  // 32'hf953441b;
    ram_cell[     244] = 32'h0;  // 32'hf490b06d;
    ram_cell[     245] = 32'h0;  // 32'h58b85a43;
    ram_cell[     246] = 32'h0;  // 32'hfbf09bb5;
    ram_cell[     247] = 32'h0;  // 32'he98f592e;
    ram_cell[     248] = 32'h0;  // 32'h48f87daa;
    ram_cell[     249] = 32'h0;  // 32'h1b9cbb7a;
    ram_cell[     250] = 32'h0;  // 32'h27436102;
    ram_cell[     251] = 32'h0;  // 32'h008e7c55;
    ram_cell[     252] = 32'h0;  // 32'hb1f4f270;
    ram_cell[     253] = 32'h0;  // 32'h8f896ac8;
    ram_cell[     254] = 32'h0;  // 32'h353e3855;
    ram_cell[     255] = 32'h0;  // 32'h2a60d344;
    // src matrix A
    ram_cell[     256] = 32'h582b69f0;
    ram_cell[     257] = 32'h51ce9689;
    ram_cell[     258] = 32'h6df60a30;
    ram_cell[     259] = 32'h31aaf4f8;
    ram_cell[     260] = 32'ha347ba15;
    ram_cell[     261] = 32'h6dddeae0;
    ram_cell[     262] = 32'hd39c4610;
    ram_cell[     263] = 32'h83713e59;
    ram_cell[     264] = 32'h93fe275d;
    ram_cell[     265] = 32'h9e105273;
    ram_cell[     266] = 32'h596529e2;
    ram_cell[     267] = 32'h594c266d;
    ram_cell[     268] = 32'ha439671e;
    ram_cell[     269] = 32'hf4c7bcb8;
    ram_cell[     270] = 32'hdbd7c55e;
    ram_cell[     271] = 32'h84734d55;
    ram_cell[     272] = 32'h19e06240;
    ram_cell[     273] = 32'h50cc0438;
    ram_cell[     274] = 32'hbcc724b0;
    ram_cell[     275] = 32'h2dbbea6a;
    ram_cell[     276] = 32'hdb12498a;
    ram_cell[     277] = 32'haeaae861;
    ram_cell[     278] = 32'h8fd340a8;
    ram_cell[     279] = 32'hc5cacfe0;
    ram_cell[     280] = 32'h03792e32;
    ram_cell[     281] = 32'he6a076ba;
    ram_cell[     282] = 32'h9f3e02e5;
    ram_cell[     283] = 32'h9f04cbef;
    ram_cell[     284] = 32'hb6e10fdb;
    ram_cell[     285] = 32'hc971e029;
    ram_cell[     286] = 32'hf85e435e;
    ram_cell[     287] = 32'h61be456a;
    ram_cell[     288] = 32'h01644492;
    ram_cell[     289] = 32'h4000a172;
    ram_cell[     290] = 32'hc86a92c8;
    ram_cell[     291] = 32'hb80bf815;
    ram_cell[     292] = 32'h1e962787;
    ram_cell[     293] = 32'h352f9f8a;
    ram_cell[     294] = 32'h86063a26;
    ram_cell[     295] = 32'h34162166;
    ram_cell[     296] = 32'h9250a5ea;
    ram_cell[     297] = 32'h27e780f2;
    ram_cell[     298] = 32'hcd048d2a;
    ram_cell[     299] = 32'h626cd2b4;
    ram_cell[     300] = 32'h284eb6dd;
    ram_cell[     301] = 32'h50e4c5f4;
    ram_cell[     302] = 32'h5089ab16;
    ram_cell[     303] = 32'hc1e92878;
    ram_cell[     304] = 32'h26c9ca00;
    ram_cell[     305] = 32'h8810bb49;
    ram_cell[     306] = 32'hee6a91cb;
    ram_cell[     307] = 32'h03159b23;
    ram_cell[     308] = 32'h06df14a7;
    ram_cell[     309] = 32'hf53a89d3;
    ram_cell[     310] = 32'h0c79fa68;
    ram_cell[     311] = 32'h727ed48b;
    ram_cell[     312] = 32'h7cc05a97;
    ram_cell[     313] = 32'hfa8c2dbd;
    ram_cell[     314] = 32'h4f36758e;
    ram_cell[     315] = 32'hd7b81a7d;
    ram_cell[     316] = 32'hd89dbd69;
    ram_cell[     317] = 32'h3ffa39b8;
    ram_cell[     318] = 32'hd2db458f;
    ram_cell[     319] = 32'h94939a03;
    ram_cell[     320] = 32'hd53786e2;
    ram_cell[     321] = 32'he4fafffc;
    ram_cell[     322] = 32'h581cb2b9;
    ram_cell[     323] = 32'hf84d6455;
    ram_cell[     324] = 32'hb8add6e4;
    ram_cell[     325] = 32'h17476541;
    ram_cell[     326] = 32'he94d52cf;
    ram_cell[     327] = 32'h60e05ddc;
    ram_cell[     328] = 32'h6f391e66;
    ram_cell[     329] = 32'h3e9d9b0f;
    ram_cell[     330] = 32'h32fe09a5;
    ram_cell[     331] = 32'h9de739c7;
    ram_cell[     332] = 32'hb31f1467;
    ram_cell[     333] = 32'h1b564c59;
    ram_cell[     334] = 32'hd4e581ec;
    ram_cell[     335] = 32'h2584afe6;
    ram_cell[     336] = 32'he5f6c41c;
    ram_cell[     337] = 32'hcaf8ec09;
    ram_cell[     338] = 32'h4c27b127;
    ram_cell[     339] = 32'h7e57e60a;
    ram_cell[     340] = 32'h1521371b;
    ram_cell[     341] = 32'hc581b713;
    ram_cell[     342] = 32'h5754957d;
    ram_cell[     343] = 32'he7c9e08b;
    ram_cell[     344] = 32'h7893ae47;
    ram_cell[     345] = 32'h3fa314a3;
    ram_cell[     346] = 32'hea726fd3;
    ram_cell[     347] = 32'h0f981161;
    ram_cell[     348] = 32'he82bf8b3;
    ram_cell[     349] = 32'heb44990f;
    ram_cell[     350] = 32'hc636902f;
    ram_cell[     351] = 32'h6636eb73;
    ram_cell[     352] = 32'hafa3256a;
    ram_cell[     353] = 32'h696b2479;
    ram_cell[     354] = 32'hbf9bfa5e;
    ram_cell[     355] = 32'h3411f2e5;
    ram_cell[     356] = 32'h8f9247b3;
    ram_cell[     357] = 32'h6c6c1f24;
    ram_cell[     358] = 32'h5794a1d2;
    ram_cell[     359] = 32'hb4d97a52;
    ram_cell[     360] = 32'hefd02767;
    ram_cell[     361] = 32'h0a0f8841;
    ram_cell[     362] = 32'h033d1476;
    ram_cell[     363] = 32'h354c6816;
    ram_cell[     364] = 32'h679b71b7;
    ram_cell[     365] = 32'hab313819;
    ram_cell[     366] = 32'h7f057f18;
    ram_cell[     367] = 32'h68bbc514;
    ram_cell[     368] = 32'h2db2063c;
    ram_cell[     369] = 32'h9ff1fce0;
    ram_cell[     370] = 32'he7a48509;
    ram_cell[     371] = 32'hb086d795;
    ram_cell[     372] = 32'h59575a37;
    ram_cell[     373] = 32'h74a299d6;
    ram_cell[     374] = 32'h88acbab4;
    ram_cell[     375] = 32'ha2c52fa7;
    ram_cell[     376] = 32'h4b5ad5aa;
    ram_cell[     377] = 32'h6271599d;
    ram_cell[     378] = 32'had9ce3b3;
    ram_cell[     379] = 32'ha742aff1;
    ram_cell[     380] = 32'hbf66c93a;
    ram_cell[     381] = 32'h06dc403a;
    ram_cell[     382] = 32'h7a84837b;
    ram_cell[     383] = 32'h0dcbad01;
    ram_cell[     384] = 32'hdfebfde6;
    ram_cell[     385] = 32'h37b5cabd;
    ram_cell[     386] = 32'h1638112d;
    ram_cell[     387] = 32'h92c87de9;
    ram_cell[     388] = 32'h2a9475ec;
    ram_cell[     389] = 32'hbddae7b4;
    ram_cell[     390] = 32'h9dd4b580;
    ram_cell[     391] = 32'h09cb51bc;
    ram_cell[     392] = 32'hf5105c94;
    ram_cell[     393] = 32'h99de9d04;
    ram_cell[     394] = 32'h7718cbea;
    ram_cell[     395] = 32'h00d17587;
    ram_cell[     396] = 32'he079e848;
    ram_cell[     397] = 32'h9fb0453e;
    ram_cell[     398] = 32'hc27961be;
    ram_cell[     399] = 32'h5274959a;
    ram_cell[     400] = 32'hb0f9c507;
    ram_cell[     401] = 32'h089f513a;
    ram_cell[     402] = 32'h9accf5d0;
    ram_cell[     403] = 32'h1ff68cc3;
    ram_cell[     404] = 32'h7d92964e;
    ram_cell[     405] = 32'h3ede9b91;
    ram_cell[     406] = 32'h67a75e6e;
    ram_cell[     407] = 32'hf5914b1d;
    ram_cell[     408] = 32'h8ad9527d;
    ram_cell[     409] = 32'hd6d888c2;
    ram_cell[     410] = 32'h9b28aefb;
    ram_cell[     411] = 32'h20d7fa02;
    ram_cell[     412] = 32'ha909989a;
    ram_cell[     413] = 32'hebe53bbb;
    ram_cell[     414] = 32'h7ff4e880;
    ram_cell[     415] = 32'h260eeeb4;
    ram_cell[     416] = 32'h54250716;
    ram_cell[     417] = 32'h38074c33;
    ram_cell[     418] = 32'hb4d09c18;
    ram_cell[     419] = 32'hcda6247f;
    ram_cell[     420] = 32'h72548b19;
    ram_cell[     421] = 32'hb51d6ad6;
    ram_cell[     422] = 32'h20f6104a;
    ram_cell[     423] = 32'h648cc9b9;
    ram_cell[     424] = 32'h9648689f;
    ram_cell[     425] = 32'h090c7c78;
    ram_cell[     426] = 32'h4f6dae9d;
    ram_cell[     427] = 32'h267e125a;
    ram_cell[     428] = 32'hf67f7418;
    ram_cell[     429] = 32'hc83718c8;
    ram_cell[     430] = 32'h5931f296;
    ram_cell[     431] = 32'h84450b4c;
    ram_cell[     432] = 32'h516c2076;
    ram_cell[     433] = 32'h8e438338;
    ram_cell[     434] = 32'he7a9b7db;
    ram_cell[     435] = 32'h8c611d89;
    ram_cell[     436] = 32'hd9c8e0b2;
    ram_cell[     437] = 32'h65f7ca74;
    ram_cell[     438] = 32'h62001329;
    ram_cell[     439] = 32'h1b093168;
    ram_cell[     440] = 32'h0de564e4;
    ram_cell[     441] = 32'h84865381;
    ram_cell[     442] = 32'hf599d618;
    ram_cell[     443] = 32'h6f6fa54a;
    ram_cell[     444] = 32'h3ab374c6;
    ram_cell[     445] = 32'h7e72050d;
    ram_cell[     446] = 32'h469bf8aa;
    ram_cell[     447] = 32'h015b6aea;
    ram_cell[     448] = 32'hbd94e873;
    ram_cell[     449] = 32'h7c20c98c;
    ram_cell[     450] = 32'h9706f109;
    ram_cell[     451] = 32'h233214b1;
    ram_cell[     452] = 32'h846d2e2a;
    ram_cell[     453] = 32'h703c551f;
    ram_cell[     454] = 32'h253b1dad;
    ram_cell[     455] = 32'h67ea62c1;
    ram_cell[     456] = 32'h31927431;
    ram_cell[     457] = 32'hb6ff9a14;
    ram_cell[     458] = 32'hf81e2c7c;
    ram_cell[     459] = 32'ha67d7339;
    ram_cell[     460] = 32'h7768d078;
    ram_cell[     461] = 32'h5289eced;
    ram_cell[     462] = 32'h8f7c16d8;
    ram_cell[     463] = 32'h18960fbf;
    ram_cell[     464] = 32'he140ee34;
    ram_cell[     465] = 32'hd562589f;
    ram_cell[     466] = 32'h74d42090;
    ram_cell[     467] = 32'ha27da205;
    ram_cell[     468] = 32'h22327bba;
    ram_cell[     469] = 32'h26ccc22f;
    ram_cell[     470] = 32'hc8cc9997;
    ram_cell[     471] = 32'h938bdb0e;
    ram_cell[     472] = 32'h5b08c90c;
    ram_cell[     473] = 32'h6da9e260;
    ram_cell[     474] = 32'h7e90d094;
    ram_cell[     475] = 32'h70ade8b0;
    ram_cell[     476] = 32'h09210207;
    ram_cell[     477] = 32'h9dfabb5c;
    ram_cell[     478] = 32'hcbbeaaf7;
    ram_cell[     479] = 32'h24855b4e;
    ram_cell[     480] = 32'hd8afcb1a;
    ram_cell[     481] = 32'h4792f8f3;
    ram_cell[     482] = 32'hb0193459;
    ram_cell[     483] = 32'ha85bb2a7;
    ram_cell[     484] = 32'he09ea0f7;
    ram_cell[     485] = 32'h90d17d06;
    ram_cell[     486] = 32'hafc8f2de;
    ram_cell[     487] = 32'h9df2d4e8;
    ram_cell[     488] = 32'h5685a816;
    ram_cell[     489] = 32'h42ba14fc;
    ram_cell[     490] = 32'h6202b37d;
    ram_cell[     491] = 32'h5ab38de1;
    ram_cell[     492] = 32'hd4ebe46e;
    ram_cell[     493] = 32'hffdba967;
    ram_cell[     494] = 32'h672b781c;
    ram_cell[     495] = 32'hae03d008;
    ram_cell[     496] = 32'h085cd778;
    ram_cell[     497] = 32'h51d87476;
    ram_cell[     498] = 32'hf9b3f08c;
    ram_cell[     499] = 32'hbd7dcbfb;
    ram_cell[     500] = 32'h6cc32203;
    ram_cell[     501] = 32'h27ae0dd1;
    ram_cell[     502] = 32'hf8207d77;
    ram_cell[     503] = 32'h8ff36f13;
    ram_cell[     504] = 32'hc4e93c8f;
    ram_cell[     505] = 32'hff8b6769;
    ram_cell[     506] = 32'h4d536513;
    ram_cell[     507] = 32'hdd984e38;
    ram_cell[     508] = 32'h7f62caed;
    ram_cell[     509] = 32'h733d9a2a;
    ram_cell[     510] = 32'h18318a10;
    ram_cell[     511] = 32'h16c8b2c6;
    // src matrix B
    ram_cell[     512] = 32'h7d0f83f4;
    ram_cell[     513] = 32'hbec2eb70;
    ram_cell[     514] = 32'hc67e34b2;
    ram_cell[     515] = 32'h9bf6a1a9;
    ram_cell[     516] = 32'h33df369e;
    ram_cell[     517] = 32'h35bc783a;
    ram_cell[     518] = 32'hbc8deb4c;
    ram_cell[     519] = 32'h209db151;
    ram_cell[     520] = 32'hcc3f8199;
    ram_cell[     521] = 32'hd03d6539;
    ram_cell[     522] = 32'hca4e661f;
    ram_cell[     523] = 32'h63e06fd1;
    ram_cell[     524] = 32'hf21e9219;
    ram_cell[     525] = 32'h320fa91d;
    ram_cell[     526] = 32'h419de37b;
    ram_cell[     527] = 32'h10294c9b;
    ram_cell[     528] = 32'h118514a2;
    ram_cell[     529] = 32'h5748d138;
    ram_cell[     530] = 32'h61f11474;
    ram_cell[     531] = 32'h35bbbb0e;
    ram_cell[     532] = 32'h16971e02;
    ram_cell[     533] = 32'hd369a6b0;
    ram_cell[     534] = 32'h823bed99;
    ram_cell[     535] = 32'h09b2ba3d;
    ram_cell[     536] = 32'h09460fb1;
    ram_cell[     537] = 32'h63ecd25c;
    ram_cell[     538] = 32'hd2c8ac18;
    ram_cell[     539] = 32'h945c87f6;
    ram_cell[     540] = 32'h1c0de22e;
    ram_cell[     541] = 32'hf54afbd1;
    ram_cell[     542] = 32'h9c223df4;
    ram_cell[     543] = 32'h9c5e30eb;
    ram_cell[     544] = 32'h0ab089e1;
    ram_cell[     545] = 32'h9757ec53;
    ram_cell[     546] = 32'h32f0f6cf;
    ram_cell[     547] = 32'hfecfaa71;
    ram_cell[     548] = 32'h57889072;
    ram_cell[     549] = 32'h169ac034;
    ram_cell[     550] = 32'h5d3cdfce;
    ram_cell[     551] = 32'hecaed177;
    ram_cell[     552] = 32'h0a7623c8;
    ram_cell[     553] = 32'hd42d9355;
    ram_cell[     554] = 32'h86aee6b4;
    ram_cell[     555] = 32'hef403b93;
    ram_cell[     556] = 32'h64c7a1af;
    ram_cell[     557] = 32'he4e44793;
    ram_cell[     558] = 32'h2ca884e4;
    ram_cell[     559] = 32'h84abab8d;
    ram_cell[     560] = 32'h0d837f3e;
    ram_cell[     561] = 32'h6ab1f0f6;
    ram_cell[     562] = 32'h1a0e5479;
    ram_cell[     563] = 32'h8ff64ae3;
    ram_cell[     564] = 32'h47a9e88e;
    ram_cell[     565] = 32'he41a01fe;
    ram_cell[     566] = 32'h071113ff;
    ram_cell[     567] = 32'hdde55a74;
    ram_cell[     568] = 32'hf22fe512;
    ram_cell[     569] = 32'h5365a9ed;
    ram_cell[     570] = 32'h6ad67a68;
    ram_cell[     571] = 32'h2d8958c8;
    ram_cell[     572] = 32'hb474d3f4;
    ram_cell[     573] = 32'hf9521bed;
    ram_cell[     574] = 32'hda33bc17;
    ram_cell[     575] = 32'heee32948;
    ram_cell[     576] = 32'h8f34f2bf;
    ram_cell[     577] = 32'hb6515857;
    ram_cell[     578] = 32'ha5abfefe;
    ram_cell[     579] = 32'hc89fec03;
    ram_cell[     580] = 32'h505090e3;
    ram_cell[     581] = 32'h6d869c0d;
    ram_cell[     582] = 32'h79415e33;
    ram_cell[     583] = 32'hd0913a83;
    ram_cell[     584] = 32'h3c188d0f;
    ram_cell[     585] = 32'h7e8ad9b5;
    ram_cell[     586] = 32'ha890567a;
    ram_cell[     587] = 32'hc9fcdba8;
    ram_cell[     588] = 32'hd7473126;
    ram_cell[     589] = 32'h563ca017;
    ram_cell[     590] = 32'hd5fad3b4;
    ram_cell[     591] = 32'h5315086b;
    ram_cell[     592] = 32'h145c7711;
    ram_cell[     593] = 32'h675ea891;
    ram_cell[     594] = 32'he7db0670;
    ram_cell[     595] = 32'h75d2b1ba;
    ram_cell[     596] = 32'h5ede696c;
    ram_cell[     597] = 32'he911c2e8;
    ram_cell[     598] = 32'h16500762;
    ram_cell[     599] = 32'he8a50708;
    ram_cell[     600] = 32'h10c19492;
    ram_cell[     601] = 32'h38b974e4;
    ram_cell[     602] = 32'h74c7f7b9;
    ram_cell[     603] = 32'h3d371b06;
    ram_cell[     604] = 32'h73c59cd9;
    ram_cell[     605] = 32'hc2f57e0e;
    ram_cell[     606] = 32'h9c37d675;
    ram_cell[     607] = 32'hb2736485;
    ram_cell[     608] = 32'haf0fe3f0;
    ram_cell[     609] = 32'h044a282c;
    ram_cell[     610] = 32'h77102b42;
    ram_cell[     611] = 32'h92acd2a4;
    ram_cell[     612] = 32'hb7f958df;
    ram_cell[     613] = 32'h9af7bd4e;
    ram_cell[     614] = 32'h1c7e2762;
    ram_cell[     615] = 32'h14b97b4b;
    ram_cell[     616] = 32'haf80ec24;
    ram_cell[     617] = 32'h4a061d25;
    ram_cell[     618] = 32'hcdcd4edf;
    ram_cell[     619] = 32'h3beb32ba;
    ram_cell[     620] = 32'ha83b5651;
    ram_cell[     621] = 32'h0ec90509;
    ram_cell[     622] = 32'hdc6bc44b;
    ram_cell[     623] = 32'h0ec5107e;
    ram_cell[     624] = 32'h67e80a20;
    ram_cell[     625] = 32'hcc2b088d;
    ram_cell[     626] = 32'hd80e8b15;
    ram_cell[     627] = 32'hf4e58d23;
    ram_cell[     628] = 32'h554781cc;
    ram_cell[     629] = 32'hfdad66ba;
    ram_cell[     630] = 32'hcae0bd15;
    ram_cell[     631] = 32'h609054f1;
    ram_cell[     632] = 32'hd7270209;
    ram_cell[     633] = 32'h17342cc1;
    ram_cell[     634] = 32'hd8b9cd1a;
    ram_cell[     635] = 32'h84cf48ee;
    ram_cell[     636] = 32'h4993ff84;
    ram_cell[     637] = 32'h1dcad038;
    ram_cell[     638] = 32'h882984ec;
    ram_cell[     639] = 32'h7f581a02;
    ram_cell[     640] = 32'hdb51a6b3;
    ram_cell[     641] = 32'h1b1e1b19;
    ram_cell[     642] = 32'h66e6d820;
    ram_cell[     643] = 32'hb98460cf;
    ram_cell[     644] = 32'h70513277;
    ram_cell[     645] = 32'h7c54e659;
    ram_cell[     646] = 32'h58a4b338;
    ram_cell[     647] = 32'he884dd4e;
    ram_cell[     648] = 32'h370ba89f;
    ram_cell[     649] = 32'h6a229fba;
    ram_cell[     650] = 32'hbd9149a5;
    ram_cell[     651] = 32'h03420759;
    ram_cell[     652] = 32'h3c8be288;
    ram_cell[     653] = 32'hb91f6f02;
    ram_cell[     654] = 32'h8a77882c;
    ram_cell[     655] = 32'hfffbc29a;
    ram_cell[     656] = 32'h3bcc8106;
    ram_cell[     657] = 32'h75fe243d;
    ram_cell[     658] = 32'hf3576913;
    ram_cell[     659] = 32'hc8f9575f;
    ram_cell[     660] = 32'ha0195ee1;
    ram_cell[     661] = 32'h10d96610;
    ram_cell[     662] = 32'h2246b2fc;
    ram_cell[     663] = 32'h9b09f00c;
    ram_cell[     664] = 32'ha1127a50;
    ram_cell[     665] = 32'hb72f3eff;
    ram_cell[     666] = 32'h0b48343c;
    ram_cell[     667] = 32'hd5e0c288;
    ram_cell[     668] = 32'h044e591a;
    ram_cell[     669] = 32'h24503a9a;
    ram_cell[     670] = 32'hfaece9ed;
    ram_cell[     671] = 32'h5319a9d2;
    ram_cell[     672] = 32'he1ff3f98;
    ram_cell[     673] = 32'h781d2eb7;
    ram_cell[     674] = 32'h947e1be3;
    ram_cell[     675] = 32'h5c2930ec;
    ram_cell[     676] = 32'h137e1c46;
    ram_cell[     677] = 32'he5d4571a;
    ram_cell[     678] = 32'h6552e592;
    ram_cell[     679] = 32'hd8880762;
    ram_cell[     680] = 32'h6efa2e45;
    ram_cell[     681] = 32'h01657408;
    ram_cell[     682] = 32'h5a009166;
    ram_cell[     683] = 32'h276d4fa2;
    ram_cell[     684] = 32'h0b355fae;
    ram_cell[     685] = 32'he96e31e6;
    ram_cell[     686] = 32'h87529425;
    ram_cell[     687] = 32'h59c6c94b;
    ram_cell[     688] = 32'h1af46c36;
    ram_cell[     689] = 32'h9700b58f;
    ram_cell[     690] = 32'h8b53d6b9;
    ram_cell[     691] = 32'h4d8527ca;
    ram_cell[     692] = 32'h6932ce62;
    ram_cell[     693] = 32'h3c493d41;
    ram_cell[     694] = 32'hbcc71b0f;
    ram_cell[     695] = 32'h925783e0;
    ram_cell[     696] = 32'hd70293f7;
    ram_cell[     697] = 32'hd321f4ce;
    ram_cell[     698] = 32'hce311965;
    ram_cell[     699] = 32'h1c440452;
    ram_cell[     700] = 32'h3b87891d;
    ram_cell[     701] = 32'h2fd5e8d5;
    ram_cell[     702] = 32'h7f39a12a;
    ram_cell[     703] = 32'h7bb8d5fd;
    ram_cell[     704] = 32'h6a9246b8;
    ram_cell[     705] = 32'h657718cd;
    ram_cell[     706] = 32'h7ab1f663;
    ram_cell[     707] = 32'he4bd04d2;
    ram_cell[     708] = 32'hd3ece95b;
    ram_cell[     709] = 32'he9432517;
    ram_cell[     710] = 32'h1d8bc922;
    ram_cell[     711] = 32'heb469cef;
    ram_cell[     712] = 32'h962077fc;
    ram_cell[     713] = 32'ha784595f;
    ram_cell[     714] = 32'hd8f47335;
    ram_cell[     715] = 32'h60c71b1a;
    ram_cell[     716] = 32'h21ea577e;
    ram_cell[     717] = 32'h9a5de6c3;
    ram_cell[     718] = 32'h5e185dc0;
    ram_cell[     719] = 32'hf943439f;
    ram_cell[     720] = 32'h3f8c5123;
    ram_cell[     721] = 32'h6c3606f7;
    ram_cell[     722] = 32'h1b1a2c93;
    ram_cell[     723] = 32'h6f6c30ff;
    ram_cell[     724] = 32'h80e1085e;
    ram_cell[     725] = 32'h693afca3;
    ram_cell[     726] = 32'h1218db31;
    ram_cell[     727] = 32'ha72a21f9;
    ram_cell[     728] = 32'h282921b5;
    ram_cell[     729] = 32'h0b7000d0;
    ram_cell[     730] = 32'h63a49d7d;
    ram_cell[     731] = 32'h45d5e0b7;
    ram_cell[     732] = 32'h2c3f54f9;
    ram_cell[     733] = 32'ha0989001;
    ram_cell[     734] = 32'h71637ecf;
    ram_cell[     735] = 32'h1550d3e6;
    ram_cell[     736] = 32'h3fe22ed2;
    ram_cell[     737] = 32'h406883e0;
    ram_cell[     738] = 32'h55cc5836;
    ram_cell[     739] = 32'h7cdd08ea;
    ram_cell[     740] = 32'h02d5c154;
    ram_cell[     741] = 32'h9d472a0a;
    ram_cell[     742] = 32'h27bc52d9;
    ram_cell[     743] = 32'h7ec42e71;
    ram_cell[     744] = 32'hfd73856a;
    ram_cell[     745] = 32'hf93b1fba;
    ram_cell[     746] = 32'hd8e9cb7a;
    ram_cell[     747] = 32'h3045adc7;
    ram_cell[     748] = 32'h4358ceff;
    ram_cell[     749] = 32'ha6ae7160;
    ram_cell[     750] = 32'h0d395dda;
    ram_cell[     751] = 32'h58af480a;
    ram_cell[     752] = 32'h91c91e2a;
    ram_cell[     753] = 32'hb9cce61d;
    ram_cell[     754] = 32'h312d05b1;
    ram_cell[     755] = 32'h7d83c69f;
    ram_cell[     756] = 32'h33abb743;
    ram_cell[     757] = 32'haeed0682;
    ram_cell[     758] = 32'h91bf6c4f;
    ram_cell[     759] = 32'hd6348bab;
    ram_cell[     760] = 32'hbed13d24;
    ram_cell[     761] = 32'h98088dfb;
    ram_cell[     762] = 32'h3047ddff;
    ram_cell[     763] = 32'h67dd97ff;
    ram_cell[     764] = 32'h0e8c2d44;
    ram_cell[     765] = 32'h9b8ffa26;
    ram_cell[     766] = 32'h6eb419c6;
    ram_cell[     767] = 32'h576a1f6e;
end

endmodule
