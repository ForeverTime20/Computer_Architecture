
module mem #(                   // 
    parameter  ADDR_LEN  = 11   // 
) (
    input  clk, rst,
    input  [ADDR_LEN-1:0] addr, // memory address
    output reg [31:0] rd_data,  // data read out
    input  wr_req,
    input  [31:0] wr_data       // data write in
);
localparam MEM_SIZE = 1<<ADDR_LEN;
reg [31:0] ram_cell [MEM_SIZE];

always @ (posedge clk or posedge rst)
    if(rst)
        rd_data <= 0;
    else
        rd_data <= ram_cell[addr];

always @ (posedge clk)
    if(wr_req) 
        ram_cell[addr] <= wr_data;

initial begin
    // dst matrix C
    ram_cell[       0] = 32'h0;  // 32'ha26db41c;
    ram_cell[       1] = 32'h0;  // 32'h74cb6ca5;
    ram_cell[       2] = 32'h0;  // 32'hff32579b;
    ram_cell[       3] = 32'h0;  // 32'hd797efa4;
    ram_cell[       4] = 32'h0;  // 32'h9bf7066f;
    ram_cell[       5] = 32'h0;  // 32'he9e3c4b6;
    ram_cell[       6] = 32'h0;  // 32'h92ced85c;
    ram_cell[       7] = 32'h0;  // 32'h366fb5b2;
    ram_cell[       8] = 32'h0;  // 32'h4d7ff636;
    ram_cell[       9] = 32'h0;  // 32'hab2c9499;
    ram_cell[      10] = 32'h0;  // 32'h4acc56bf;
    ram_cell[      11] = 32'h0;  // 32'haa47c206;
    ram_cell[      12] = 32'h0;  // 32'h944553dc;
    ram_cell[      13] = 32'h0;  // 32'h6214845a;
    ram_cell[      14] = 32'h0;  // 32'h9a470127;
    ram_cell[      15] = 32'h0;  // 32'h3717f0d8;
    ram_cell[      16] = 32'h0;  // 32'hf45f6ad1;
    ram_cell[      17] = 32'h0;  // 32'h59a3f79f;
    ram_cell[      18] = 32'h0;  // 32'hef3b93cc;
    ram_cell[      19] = 32'h0;  // 32'hee0661a7;
    ram_cell[      20] = 32'h0;  // 32'haed9bcaa;
    ram_cell[      21] = 32'h0;  // 32'h75cfddff;
    ram_cell[      22] = 32'h0;  // 32'h23f8270f;
    ram_cell[      23] = 32'h0;  // 32'h1c7fa4bb;
    ram_cell[      24] = 32'h0;  // 32'hac913e2d;
    ram_cell[      25] = 32'h0;  // 32'h1bc52a1a;
    ram_cell[      26] = 32'h0;  // 32'h4c2b4641;
    ram_cell[      27] = 32'h0;  // 32'h690a780d;
    ram_cell[      28] = 32'h0;  // 32'h19d17071;
    ram_cell[      29] = 32'h0;  // 32'h9361a787;
    ram_cell[      30] = 32'h0;  // 32'h9a9cb213;
    ram_cell[      31] = 32'h0;  // 32'h7f3a5f16;
    ram_cell[      32] = 32'h0;  // 32'hb38edc4d;
    ram_cell[      33] = 32'h0;  // 32'h835af690;
    ram_cell[      34] = 32'h0;  // 32'h5dade76b;
    ram_cell[      35] = 32'h0;  // 32'hb0b7d5de;
    ram_cell[      36] = 32'h0;  // 32'h18e3662a;
    ram_cell[      37] = 32'h0;  // 32'h82f85fac;
    ram_cell[      38] = 32'h0;  // 32'h4730c548;
    ram_cell[      39] = 32'h0;  // 32'h5c7e8403;
    ram_cell[      40] = 32'h0;  // 32'h53b91fd0;
    ram_cell[      41] = 32'h0;  // 32'hc8c47689;
    ram_cell[      42] = 32'h0;  // 32'hf88cfffa;
    ram_cell[      43] = 32'h0;  // 32'hfea2e714;
    ram_cell[      44] = 32'h0;  // 32'hb4a12317;
    ram_cell[      45] = 32'h0;  // 32'h4ff933e5;
    ram_cell[      46] = 32'h0;  // 32'hba2627f9;
    ram_cell[      47] = 32'h0;  // 32'h8d625462;
    ram_cell[      48] = 32'h0;  // 32'h245e7e8b;
    ram_cell[      49] = 32'h0;  // 32'hc06dc7ff;
    ram_cell[      50] = 32'h0;  // 32'h91dccd7f;
    ram_cell[      51] = 32'h0;  // 32'h8595b782;
    ram_cell[      52] = 32'h0;  // 32'hc207f873;
    ram_cell[      53] = 32'h0;  // 32'h769ed49e;
    ram_cell[      54] = 32'h0;  // 32'hd987a1d6;
    ram_cell[      55] = 32'h0;  // 32'ha03e0cef;
    ram_cell[      56] = 32'h0;  // 32'h48e7c9a3;
    ram_cell[      57] = 32'h0;  // 32'h4809e56f;
    ram_cell[      58] = 32'h0;  // 32'h865e7830;
    ram_cell[      59] = 32'h0;  // 32'h036ccb6f;
    ram_cell[      60] = 32'h0;  // 32'h20edf680;
    ram_cell[      61] = 32'h0;  // 32'hf3bb56a3;
    ram_cell[      62] = 32'h0;  // 32'hbb0942d2;
    ram_cell[      63] = 32'h0;  // 32'hfe793901;
    ram_cell[      64] = 32'h0;  // 32'hf8247682;
    ram_cell[      65] = 32'h0;  // 32'h21123125;
    ram_cell[      66] = 32'h0;  // 32'h25edbd64;
    ram_cell[      67] = 32'h0;  // 32'hdb1b8863;
    ram_cell[      68] = 32'h0;  // 32'hc46ff5c9;
    ram_cell[      69] = 32'h0;  // 32'hfc536859;
    ram_cell[      70] = 32'h0;  // 32'h48ed6694;
    ram_cell[      71] = 32'h0;  // 32'h90c0fa33;
    ram_cell[      72] = 32'h0;  // 32'h50bbf697;
    ram_cell[      73] = 32'h0;  // 32'h8945e649;
    ram_cell[      74] = 32'h0;  // 32'h544f626e;
    ram_cell[      75] = 32'h0;  // 32'he2e5df07;
    ram_cell[      76] = 32'h0;  // 32'hf8824c4c;
    ram_cell[      77] = 32'h0;  // 32'h93c9e402;
    ram_cell[      78] = 32'h0;  // 32'h12c5fc19;
    ram_cell[      79] = 32'h0;  // 32'h9f6ca5d3;
    ram_cell[      80] = 32'h0;  // 32'h0b7389ba;
    ram_cell[      81] = 32'h0;  // 32'h36d12173;
    ram_cell[      82] = 32'h0;  // 32'h326ca586;
    ram_cell[      83] = 32'h0;  // 32'hf717a06b;
    ram_cell[      84] = 32'h0;  // 32'h3064c7bd;
    ram_cell[      85] = 32'h0;  // 32'hd0c6d090;
    ram_cell[      86] = 32'h0;  // 32'h6e0f7f44;
    ram_cell[      87] = 32'h0;  // 32'h81fb4f83;
    ram_cell[      88] = 32'h0;  // 32'h9f121e47;
    ram_cell[      89] = 32'h0;  // 32'h57e950a6;
    ram_cell[      90] = 32'h0;  // 32'h8d59c673;
    ram_cell[      91] = 32'h0;  // 32'hd1ccd403;
    ram_cell[      92] = 32'h0;  // 32'hacb4afcb;
    ram_cell[      93] = 32'h0;  // 32'h3d1c6482;
    ram_cell[      94] = 32'h0;  // 32'h0249869f;
    ram_cell[      95] = 32'h0;  // 32'h4cfdf2e4;
    ram_cell[      96] = 32'h0;  // 32'h461e3e47;
    ram_cell[      97] = 32'h0;  // 32'h14392e97;
    ram_cell[      98] = 32'h0;  // 32'h36513062;
    ram_cell[      99] = 32'h0;  // 32'h7ba50c60;
    ram_cell[     100] = 32'h0;  // 32'hb3ec0cbb;
    ram_cell[     101] = 32'h0;  // 32'h120dfc4c;
    ram_cell[     102] = 32'h0;  // 32'h4ec86c93;
    ram_cell[     103] = 32'h0;  // 32'hc7282dd1;
    ram_cell[     104] = 32'h0;  // 32'h22eba432;
    ram_cell[     105] = 32'h0;  // 32'hcedff889;
    ram_cell[     106] = 32'h0;  // 32'h725a0911;
    ram_cell[     107] = 32'h0;  // 32'h1dfe5247;
    ram_cell[     108] = 32'h0;  // 32'h61acf7db;
    ram_cell[     109] = 32'h0;  // 32'h9c269701;
    ram_cell[     110] = 32'h0;  // 32'h9a059cfd;
    ram_cell[     111] = 32'h0;  // 32'hab8d490a;
    ram_cell[     112] = 32'h0;  // 32'h60a264fd;
    ram_cell[     113] = 32'h0;  // 32'hae8bd0c5;
    ram_cell[     114] = 32'h0;  // 32'h2b05dca6;
    ram_cell[     115] = 32'h0;  // 32'hb844e57a;
    ram_cell[     116] = 32'h0;  // 32'hf1dea696;
    ram_cell[     117] = 32'h0;  // 32'hfa040479;
    ram_cell[     118] = 32'h0;  // 32'h064c33c4;
    ram_cell[     119] = 32'h0;  // 32'h8a13fe1d;
    ram_cell[     120] = 32'h0;  // 32'ha7a577ba;
    ram_cell[     121] = 32'h0;  // 32'hde4b672d;
    ram_cell[     122] = 32'h0;  // 32'hccf1913e;
    ram_cell[     123] = 32'h0;  // 32'h2c95892c;
    ram_cell[     124] = 32'h0;  // 32'hb9d2faa9;
    ram_cell[     125] = 32'h0;  // 32'h9c9bd014;
    ram_cell[     126] = 32'h0;  // 32'h4adde9da;
    ram_cell[     127] = 32'h0;  // 32'hbd19ec42;
    ram_cell[     128] = 32'h0;  // 32'h30a860ef;
    ram_cell[     129] = 32'h0;  // 32'h974cd8ba;
    ram_cell[     130] = 32'h0;  // 32'h43ed9b32;
    ram_cell[     131] = 32'h0;  // 32'h1e644853;
    ram_cell[     132] = 32'h0;  // 32'h5d260b58;
    ram_cell[     133] = 32'h0;  // 32'h18354da0;
    ram_cell[     134] = 32'h0;  // 32'h29b6d164;
    ram_cell[     135] = 32'h0;  // 32'h294c44dd;
    ram_cell[     136] = 32'h0;  // 32'he19706b8;
    ram_cell[     137] = 32'h0;  // 32'h7a699426;
    ram_cell[     138] = 32'h0;  // 32'h05a82f65;
    ram_cell[     139] = 32'h0;  // 32'hdcb1fd53;
    ram_cell[     140] = 32'h0;  // 32'ha284ac03;
    ram_cell[     141] = 32'h0;  // 32'h8dad33bd;
    ram_cell[     142] = 32'h0;  // 32'h370a5534;
    ram_cell[     143] = 32'h0;  // 32'haa5bb5e9;
    ram_cell[     144] = 32'h0;  // 32'h240ea696;
    ram_cell[     145] = 32'h0;  // 32'h0b470748;
    ram_cell[     146] = 32'h0;  // 32'ha0654801;
    ram_cell[     147] = 32'h0;  // 32'h6820a261;
    ram_cell[     148] = 32'h0;  // 32'hac725d97;
    ram_cell[     149] = 32'h0;  // 32'ha790879c;
    ram_cell[     150] = 32'h0;  // 32'h47cc318f;
    ram_cell[     151] = 32'h0;  // 32'h70c848cb;
    ram_cell[     152] = 32'h0;  // 32'h9599e42e;
    ram_cell[     153] = 32'h0;  // 32'h102b3670;
    ram_cell[     154] = 32'h0;  // 32'ha4877217;
    ram_cell[     155] = 32'h0;  // 32'h0e923967;
    ram_cell[     156] = 32'h0;  // 32'h0dfaae14;
    ram_cell[     157] = 32'h0;  // 32'hf578cbe6;
    ram_cell[     158] = 32'h0;  // 32'h4c3435f2;
    ram_cell[     159] = 32'h0;  // 32'he37d8449;
    ram_cell[     160] = 32'h0;  // 32'h3d34a5ac;
    ram_cell[     161] = 32'h0;  // 32'h74381b3a;
    ram_cell[     162] = 32'h0;  // 32'h836f2049;
    ram_cell[     163] = 32'h0;  // 32'hf3a8e741;
    ram_cell[     164] = 32'h0;  // 32'h27800e8f;
    ram_cell[     165] = 32'h0;  // 32'hcd3dd97f;
    ram_cell[     166] = 32'h0;  // 32'h57661d98;
    ram_cell[     167] = 32'h0;  // 32'h8b745eb2;
    ram_cell[     168] = 32'h0;  // 32'hde1c9cc9;
    ram_cell[     169] = 32'h0;  // 32'hd500203e;
    ram_cell[     170] = 32'h0;  // 32'h4e739cb3;
    ram_cell[     171] = 32'h0;  // 32'h47c5f38b;
    ram_cell[     172] = 32'h0;  // 32'hf4142959;
    ram_cell[     173] = 32'h0;  // 32'h650c20b7;
    ram_cell[     174] = 32'h0;  // 32'h68152680;
    ram_cell[     175] = 32'h0;  // 32'hf13729ba;
    ram_cell[     176] = 32'h0;  // 32'h76219c7c;
    ram_cell[     177] = 32'h0;  // 32'h0ccaafb5;
    ram_cell[     178] = 32'h0;  // 32'h0ea0bdc9;
    ram_cell[     179] = 32'h0;  // 32'h4dd0b02c;
    ram_cell[     180] = 32'h0;  // 32'hd1ff615b;
    ram_cell[     181] = 32'h0;  // 32'h5dce0b27;
    ram_cell[     182] = 32'h0;  // 32'h84f90c9d;
    ram_cell[     183] = 32'h0;  // 32'h86f8374d;
    ram_cell[     184] = 32'h0;  // 32'h9b0e8252;
    ram_cell[     185] = 32'h0;  // 32'hc76045b3;
    ram_cell[     186] = 32'h0;  // 32'hbb2b22d5;
    ram_cell[     187] = 32'h0;  // 32'hf1c3140a;
    ram_cell[     188] = 32'h0;  // 32'h2d37e089;
    ram_cell[     189] = 32'h0;  // 32'hb98d4c71;
    ram_cell[     190] = 32'h0;  // 32'h95b643cc;
    ram_cell[     191] = 32'h0;  // 32'h35520f37;
    ram_cell[     192] = 32'h0;  // 32'hc0f83970;
    ram_cell[     193] = 32'h0;  // 32'ha6d42239;
    ram_cell[     194] = 32'h0;  // 32'hbe8781e6;
    ram_cell[     195] = 32'h0;  // 32'h4d286710;
    ram_cell[     196] = 32'h0;  // 32'h0b367605;
    ram_cell[     197] = 32'h0;  // 32'h0596f9a0;
    ram_cell[     198] = 32'h0;  // 32'he1483b58;
    ram_cell[     199] = 32'h0;  // 32'h7a964256;
    ram_cell[     200] = 32'h0;  // 32'h69f53d0b;
    ram_cell[     201] = 32'h0;  // 32'h5818aa11;
    ram_cell[     202] = 32'h0;  // 32'h6df069d1;
    ram_cell[     203] = 32'h0;  // 32'h61d94ecf;
    ram_cell[     204] = 32'h0;  // 32'hfc05a971;
    ram_cell[     205] = 32'h0;  // 32'hb65e9cea;
    ram_cell[     206] = 32'h0;  // 32'h87f41dd2;
    ram_cell[     207] = 32'h0;  // 32'h6eb51416;
    ram_cell[     208] = 32'h0;  // 32'h706c1501;
    ram_cell[     209] = 32'h0;  // 32'h20547ae9;
    ram_cell[     210] = 32'h0;  // 32'hfc22421c;
    ram_cell[     211] = 32'h0;  // 32'h27feef7b;
    ram_cell[     212] = 32'h0;  // 32'h4127bf5e;
    ram_cell[     213] = 32'h0;  // 32'hb35f2e88;
    ram_cell[     214] = 32'h0;  // 32'hea7bdd6e;
    ram_cell[     215] = 32'h0;  // 32'h9712353e;
    ram_cell[     216] = 32'h0;  // 32'hb1799290;
    ram_cell[     217] = 32'h0;  // 32'h0c190828;
    ram_cell[     218] = 32'h0;  // 32'h3a9ffef9;
    ram_cell[     219] = 32'h0;  // 32'ha3f941c0;
    ram_cell[     220] = 32'h0;  // 32'hb7a2d7d5;
    ram_cell[     221] = 32'h0;  // 32'he7fbb598;
    ram_cell[     222] = 32'h0;  // 32'h67f6f417;
    ram_cell[     223] = 32'h0;  // 32'h6afd4e56;
    ram_cell[     224] = 32'h0;  // 32'h68c7b0d0;
    ram_cell[     225] = 32'h0;  // 32'h36841ee3;
    ram_cell[     226] = 32'h0;  // 32'h0c0fdd17;
    ram_cell[     227] = 32'h0;  // 32'hce71f6e2;
    ram_cell[     228] = 32'h0;  // 32'hb3010e56;
    ram_cell[     229] = 32'h0;  // 32'hc6bd6a27;
    ram_cell[     230] = 32'h0;  // 32'h1572293f;
    ram_cell[     231] = 32'h0;  // 32'hd419445a;
    ram_cell[     232] = 32'h0;  // 32'haabc9217;
    ram_cell[     233] = 32'h0;  // 32'h84c39467;
    ram_cell[     234] = 32'h0;  // 32'h2cdd76a1;
    ram_cell[     235] = 32'h0;  // 32'h9c0d50c9;
    ram_cell[     236] = 32'h0;  // 32'h0d0f470c;
    ram_cell[     237] = 32'h0;  // 32'h0bcffcc2;
    ram_cell[     238] = 32'h0;  // 32'h55b07c94;
    ram_cell[     239] = 32'h0;  // 32'h9739a644;
    ram_cell[     240] = 32'h0;  // 32'h457b7d72;
    ram_cell[     241] = 32'h0;  // 32'hcbafcd61;
    ram_cell[     242] = 32'h0;  // 32'h023a44a7;
    ram_cell[     243] = 32'h0;  // 32'h76031a6c;
    ram_cell[     244] = 32'h0;  // 32'hc44fc99f;
    ram_cell[     245] = 32'h0;  // 32'hb989a2f1;
    ram_cell[     246] = 32'h0;  // 32'h0b43ef73;
    ram_cell[     247] = 32'h0;  // 32'h40d7828c;
    ram_cell[     248] = 32'h0;  // 32'h7edfda3a;
    ram_cell[     249] = 32'h0;  // 32'h32d6fdea;
    ram_cell[     250] = 32'h0;  // 32'hcf0e8939;
    ram_cell[     251] = 32'h0;  // 32'h252cfab2;
    ram_cell[     252] = 32'h0;  // 32'hcb356510;
    ram_cell[     253] = 32'h0;  // 32'hb948131f;
    ram_cell[     254] = 32'h0;  // 32'h6437b38b;
    ram_cell[     255] = 32'h0;  // 32'h599ad247;
    // src matrix A
    ram_cell[     256] = 32'h1fe94454;
    ram_cell[     257] = 32'h6aae6850;
    ram_cell[     258] = 32'h65a1d8e6;
    ram_cell[     259] = 32'hd9482182;
    ram_cell[     260] = 32'h1057893a;
    ram_cell[     261] = 32'h1bff2b73;
    ram_cell[     262] = 32'h7208e7a8;
    ram_cell[     263] = 32'h4824a04b;
    ram_cell[     264] = 32'haf65fca2;
    ram_cell[     265] = 32'h5c70f544;
    ram_cell[     266] = 32'hdbaa4300;
    ram_cell[     267] = 32'he14b31e3;
    ram_cell[     268] = 32'had273e0d;
    ram_cell[     269] = 32'hef31d085;
    ram_cell[     270] = 32'h240d33ff;
    ram_cell[     271] = 32'he4630e50;
    ram_cell[     272] = 32'hd5aaf86e;
    ram_cell[     273] = 32'hc6329374;
    ram_cell[     274] = 32'h3cafbd0a;
    ram_cell[     275] = 32'hbea6165b;
    ram_cell[     276] = 32'h28d45d46;
    ram_cell[     277] = 32'h03bdd3be;
    ram_cell[     278] = 32'h31f3a3d9;
    ram_cell[     279] = 32'hc09bd72f;
    ram_cell[     280] = 32'hbf2c65a3;
    ram_cell[     281] = 32'h6bdbcbd4;
    ram_cell[     282] = 32'h94fa4671;
    ram_cell[     283] = 32'h8e5c618d;
    ram_cell[     284] = 32'h31ed5fb1;
    ram_cell[     285] = 32'hb5f9c5ec;
    ram_cell[     286] = 32'h1e961a75;
    ram_cell[     287] = 32'hf697f47f;
    ram_cell[     288] = 32'h95f66c47;
    ram_cell[     289] = 32'h973696d6;
    ram_cell[     290] = 32'h0b733176;
    ram_cell[     291] = 32'hd5f9adc4;
    ram_cell[     292] = 32'h36dfe0db;
    ram_cell[     293] = 32'h0709ac1b;
    ram_cell[     294] = 32'hb91fc369;
    ram_cell[     295] = 32'h38e6d575;
    ram_cell[     296] = 32'he397047e;
    ram_cell[     297] = 32'h8848a015;
    ram_cell[     298] = 32'ha83b7520;
    ram_cell[     299] = 32'hae3b338d;
    ram_cell[     300] = 32'hd620c7ae;
    ram_cell[     301] = 32'he0bbc414;
    ram_cell[     302] = 32'he37b82c2;
    ram_cell[     303] = 32'ha023eb4c;
    ram_cell[     304] = 32'hd444def3;
    ram_cell[     305] = 32'h56778f1b;
    ram_cell[     306] = 32'hfbab8589;
    ram_cell[     307] = 32'hc9b21f33;
    ram_cell[     308] = 32'hb2a9b6aa;
    ram_cell[     309] = 32'ha9059708;
    ram_cell[     310] = 32'h914a9ec4;
    ram_cell[     311] = 32'h08ffc93d;
    ram_cell[     312] = 32'hde2349f7;
    ram_cell[     313] = 32'h92b0e43b;
    ram_cell[     314] = 32'he4b1809b;
    ram_cell[     315] = 32'ha3b4eaa0;
    ram_cell[     316] = 32'hdcb7688c;
    ram_cell[     317] = 32'h821f1589;
    ram_cell[     318] = 32'h0a0684ae;
    ram_cell[     319] = 32'h30ec036b;
    ram_cell[     320] = 32'h933bd3d6;
    ram_cell[     321] = 32'h89208cf3;
    ram_cell[     322] = 32'h1b368c75;
    ram_cell[     323] = 32'hfbf8ea82;
    ram_cell[     324] = 32'hb91665b4;
    ram_cell[     325] = 32'h841b6ea2;
    ram_cell[     326] = 32'h790c7060;
    ram_cell[     327] = 32'h13285df6;
    ram_cell[     328] = 32'h0e2e0244;
    ram_cell[     329] = 32'h01be4441;
    ram_cell[     330] = 32'h481299ed;
    ram_cell[     331] = 32'hb43ce348;
    ram_cell[     332] = 32'h3a5ae63d;
    ram_cell[     333] = 32'h5cbcd051;
    ram_cell[     334] = 32'hcbfa1362;
    ram_cell[     335] = 32'hff45b209;
    ram_cell[     336] = 32'hab8bd909;
    ram_cell[     337] = 32'h85c1e768;
    ram_cell[     338] = 32'h73b6acec;
    ram_cell[     339] = 32'h80ca13cd;
    ram_cell[     340] = 32'hf77d37b9;
    ram_cell[     341] = 32'hcc6decc7;
    ram_cell[     342] = 32'ha00fec0a;
    ram_cell[     343] = 32'h76f9f4e2;
    ram_cell[     344] = 32'h96139872;
    ram_cell[     345] = 32'hdac99847;
    ram_cell[     346] = 32'h9e0ca854;
    ram_cell[     347] = 32'h8c004d30;
    ram_cell[     348] = 32'h88aed2bb;
    ram_cell[     349] = 32'hf219cfae;
    ram_cell[     350] = 32'h53db748e;
    ram_cell[     351] = 32'hbd89be58;
    ram_cell[     352] = 32'he5ad7f0a;
    ram_cell[     353] = 32'h435f0e5d;
    ram_cell[     354] = 32'h18816d14;
    ram_cell[     355] = 32'h75299a31;
    ram_cell[     356] = 32'hf22980e2;
    ram_cell[     357] = 32'h716b1ca8;
    ram_cell[     358] = 32'h2342db41;
    ram_cell[     359] = 32'hc3c294a7;
    ram_cell[     360] = 32'h5aae14cd;
    ram_cell[     361] = 32'h2434d896;
    ram_cell[     362] = 32'haf549800;
    ram_cell[     363] = 32'hbf0e7c1e;
    ram_cell[     364] = 32'h836a6ff6;
    ram_cell[     365] = 32'h6dd3c2f9;
    ram_cell[     366] = 32'h6659e746;
    ram_cell[     367] = 32'h7acbcffc;
    ram_cell[     368] = 32'hbabae54c;
    ram_cell[     369] = 32'h8d8084ef;
    ram_cell[     370] = 32'hcc167f36;
    ram_cell[     371] = 32'h2d02260f;
    ram_cell[     372] = 32'h0e229417;
    ram_cell[     373] = 32'ha30bbe35;
    ram_cell[     374] = 32'ha754dc86;
    ram_cell[     375] = 32'h521d54ea;
    ram_cell[     376] = 32'h3de5cf23;
    ram_cell[     377] = 32'h610b8378;
    ram_cell[     378] = 32'hfc55fba1;
    ram_cell[     379] = 32'hab969078;
    ram_cell[     380] = 32'hf82e30b1;
    ram_cell[     381] = 32'h5b1cf22c;
    ram_cell[     382] = 32'hd8920c31;
    ram_cell[     383] = 32'h3edbf450;
    ram_cell[     384] = 32'h69204826;
    ram_cell[     385] = 32'h2ac0f37b;
    ram_cell[     386] = 32'h96e587df;
    ram_cell[     387] = 32'h17435b1f;
    ram_cell[     388] = 32'h60d20015;
    ram_cell[     389] = 32'h21e61a17;
    ram_cell[     390] = 32'hf0db0a70;
    ram_cell[     391] = 32'ha7e7c679;
    ram_cell[     392] = 32'hd8ab0ce1;
    ram_cell[     393] = 32'h0580115b;
    ram_cell[     394] = 32'h5acf6334;
    ram_cell[     395] = 32'h882e73a2;
    ram_cell[     396] = 32'hfe596692;
    ram_cell[     397] = 32'h4cfbb735;
    ram_cell[     398] = 32'hcb5da0d3;
    ram_cell[     399] = 32'h3b90a143;
    ram_cell[     400] = 32'h5b7bfbfb;
    ram_cell[     401] = 32'hdfb9056d;
    ram_cell[     402] = 32'h52c9af88;
    ram_cell[     403] = 32'hf852f221;
    ram_cell[     404] = 32'h39d8add5;
    ram_cell[     405] = 32'h09158939;
    ram_cell[     406] = 32'h1e629e55;
    ram_cell[     407] = 32'h426051bd;
    ram_cell[     408] = 32'hfd72b346;
    ram_cell[     409] = 32'h526e0a4e;
    ram_cell[     410] = 32'h13055142;
    ram_cell[     411] = 32'hc7d7eb92;
    ram_cell[     412] = 32'had42c995;
    ram_cell[     413] = 32'hfb581403;
    ram_cell[     414] = 32'hec975707;
    ram_cell[     415] = 32'h7fa2f0b3;
    ram_cell[     416] = 32'hfbb539e9;
    ram_cell[     417] = 32'h978c1d6d;
    ram_cell[     418] = 32'hf21b7c89;
    ram_cell[     419] = 32'hdf6070e1;
    ram_cell[     420] = 32'h20c9b5b1;
    ram_cell[     421] = 32'h25a671c3;
    ram_cell[     422] = 32'h38962b8e;
    ram_cell[     423] = 32'h7caa28cc;
    ram_cell[     424] = 32'h2512e73e;
    ram_cell[     425] = 32'h22d69b8f;
    ram_cell[     426] = 32'he137ef9d;
    ram_cell[     427] = 32'h75b001c6;
    ram_cell[     428] = 32'h2902f6f8;
    ram_cell[     429] = 32'hb367f48f;
    ram_cell[     430] = 32'h6510acbc;
    ram_cell[     431] = 32'h23db5d67;
    ram_cell[     432] = 32'h20170410;
    ram_cell[     433] = 32'hc9f4f162;
    ram_cell[     434] = 32'h29e176a5;
    ram_cell[     435] = 32'h3ee12575;
    ram_cell[     436] = 32'h2a6f7697;
    ram_cell[     437] = 32'h20c77f22;
    ram_cell[     438] = 32'hd779350f;
    ram_cell[     439] = 32'h1d391244;
    ram_cell[     440] = 32'h4bf3d23c;
    ram_cell[     441] = 32'h68dad06e;
    ram_cell[     442] = 32'hf32745d1;
    ram_cell[     443] = 32'h7324402a;
    ram_cell[     444] = 32'h42e2aa11;
    ram_cell[     445] = 32'h9517a34d;
    ram_cell[     446] = 32'h252fc187;
    ram_cell[     447] = 32'h249e6834;
    ram_cell[     448] = 32'h1bc62cf0;
    ram_cell[     449] = 32'h2e4f82fc;
    ram_cell[     450] = 32'hf2360f65;
    ram_cell[     451] = 32'hf542c1f9;
    ram_cell[     452] = 32'h138028ba;
    ram_cell[     453] = 32'h4e2d81c4;
    ram_cell[     454] = 32'h82b1a620;
    ram_cell[     455] = 32'ha8d01bb7;
    ram_cell[     456] = 32'h6a09e86b;
    ram_cell[     457] = 32'h209abede;
    ram_cell[     458] = 32'haa489129;
    ram_cell[     459] = 32'h7507fe28;
    ram_cell[     460] = 32'h01924011;
    ram_cell[     461] = 32'h8eb8e7b6;
    ram_cell[     462] = 32'h167130ed;
    ram_cell[     463] = 32'h4995408c;
    ram_cell[     464] = 32'heac777ac;
    ram_cell[     465] = 32'h3ce9e4fb;
    ram_cell[     466] = 32'ha8d44059;
    ram_cell[     467] = 32'h2a5ae8ea;
    ram_cell[     468] = 32'h5a005b9d;
    ram_cell[     469] = 32'hb926506d;
    ram_cell[     470] = 32'h4193679c;
    ram_cell[     471] = 32'hf999a9c5;
    ram_cell[     472] = 32'h05ecb53a;
    ram_cell[     473] = 32'hda09349b;
    ram_cell[     474] = 32'h817a7798;
    ram_cell[     475] = 32'h01828327;
    ram_cell[     476] = 32'h93df9d7b;
    ram_cell[     477] = 32'h56e28b36;
    ram_cell[     478] = 32'hee7bef92;
    ram_cell[     479] = 32'hb8251fa4;
    ram_cell[     480] = 32'h602f7fdb;
    ram_cell[     481] = 32'h470552bf;
    ram_cell[     482] = 32'hf153a0cc;
    ram_cell[     483] = 32'h295a6e0a;
    ram_cell[     484] = 32'habe1959a;
    ram_cell[     485] = 32'h31b4f83e;
    ram_cell[     486] = 32'hc8990de7;
    ram_cell[     487] = 32'hd41bbee1;
    ram_cell[     488] = 32'h0e4b8c28;
    ram_cell[     489] = 32'h9a6a8fa8;
    ram_cell[     490] = 32'h4554469b;
    ram_cell[     491] = 32'h54ddf730;
    ram_cell[     492] = 32'h79aae191;
    ram_cell[     493] = 32'h2a4d7750;
    ram_cell[     494] = 32'h9e25ce92;
    ram_cell[     495] = 32'h8d202931;
    ram_cell[     496] = 32'h06d9b8d7;
    ram_cell[     497] = 32'h97fa8427;
    ram_cell[     498] = 32'hcbe17bae;
    ram_cell[     499] = 32'hb6982709;
    ram_cell[     500] = 32'hd51727ec;
    ram_cell[     501] = 32'h412f73f9;
    ram_cell[     502] = 32'hcbc78393;
    ram_cell[     503] = 32'hb7ae0d62;
    ram_cell[     504] = 32'hed1afd9d;
    ram_cell[     505] = 32'had28161c;
    ram_cell[     506] = 32'heff820d9;
    ram_cell[     507] = 32'h99294d62;
    ram_cell[     508] = 32'hac4d3e31;
    ram_cell[     509] = 32'h215e2f8e;
    ram_cell[     510] = 32'hb118e94c;
    ram_cell[     511] = 32'h9de0adf1;
    // src matrix B
    ram_cell[     512] = 32'h140ca57d;
    ram_cell[     513] = 32'hb295a660;
    ram_cell[     514] = 32'h8cb0a33c;
    ram_cell[     515] = 32'h85f8f6b3;
    ram_cell[     516] = 32'h7931cdc3;
    ram_cell[     517] = 32'hce3ab3a2;
    ram_cell[     518] = 32'h015a3937;
    ram_cell[     519] = 32'ha71fa2dd;
    ram_cell[     520] = 32'h44c46369;
    ram_cell[     521] = 32'ha7260808;
    ram_cell[     522] = 32'hf6b86cbc;
    ram_cell[     523] = 32'he2eebe1f;
    ram_cell[     524] = 32'ha0a4df6d;
    ram_cell[     525] = 32'h2eb8ef40;
    ram_cell[     526] = 32'hfd485659;
    ram_cell[     527] = 32'he5dd8b70;
    ram_cell[     528] = 32'h3569407a;
    ram_cell[     529] = 32'he288dd78;
    ram_cell[     530] = 32'hffc37473;
    ram_cell[     531] = 32'hdcd590d1;
    ram_cell[     532] = 32'he99053e2;
    ram_cell[     533] = 32'h5a4d1bd0;
    ram_cell[     534] = 32'hee86f356;
    ram_cell[     535] = 32'h83d787f1;
    ram_cell[     536] = 32'h106bdd4e;
    ram_cell[     537] = 32'hfe957159;
    ram_cell[     538] = 32'h5b82badc;
    ram_cell[     539] = 32'hbbb71acd;
    ram_cell[     540] = 32'hb02a471a;
    ram_cell[     541] = 32'h700a8a89;
    ram_cell[     542] = 32'h2edcc4bc;
    ram_cell[     543] = 32'h8a9920d1;
    ram_cell[     544] = 32'h785ad3bb;
    ram_cell[     545] = 32'h784f2c36;
    ram_cell[     546] = 32'h11c8189f;
    ram_cell[     547] = 32'hb11ad439;
    ram_cell[     548] = 32'h018dcfa1;
    ram_cell[     549] = 32'h9863eb1e;
    ram_cell[     550] = 32'h0a1ea803;
    ram_cell[     551] = 32'hab6f6d1b;
    ram_cell[     552] = 32'h22e7e2ca;
    ram_cell[     553] = 32'h4cd20c97;
    ram_cell[     554] = 32'hd0c92ced;
    ram_cell[     555] = 32'he2492d6e;
    ram_cell[     556] = 32'h11eecee8;
    ram_cell[     557] = 32'hbd1ac4fd;
    ram_cell[     558] = 32'he40c624a;
    ram_cell[     559] = 32'hc29f6e2a;
    ram_cell[     560] = 32'h778b24ea;
    ram_cell[     561] = 32'h87fdddca;
    ram_cell[     562] = 32'hd2855928;
    ram_cell[     563] = 32'ha4408e7a;
    ram_cell[     564] = 32'hf766011d;
    ram_cell[     565] = 32'hf4cedf5e;
    ram_cell[     566] = 32'hb0a7e815;
    ram_cell[     567] = 32'hde25d59d;
    ram_cell[     568] = 32'h743b34a1;
    ram_cell[     569] = 32'hc2bd54ad;
    ram_cell[     570] = 32'h04055486;
    ram_cell[     571] = 32'h677a0bd4;
    ram_cell[     572] = 32'hf89a9861;
    ram_cell[     573] = 32'h4334b106;
    ram_cell[     574] = 32'hc90b5357;
    ram_cell[     575] = 32'h2d4bf52d;
    ram_cell[     576] = 32'hd39523bb;
    ram_cell[     577] = 32'h350986f9;
    ram_cell[     578] = 32'hdeeb9608;
    ram_cell[     579] = 32'he3e56a37;
    ram_cell[     580] = 32'h954ffe46;
    ram_cell[     581] = 32'h39a61d6f;
    ram_cell[     582] = 32'h87c1a265;
    ram_cell[     583] = 32'hbb800550;
    ram_cell[     584] = 32'h7d8c5998;
    ram_cell[     585] = 32'h1a12616f;
    ram_cell[     586] = 32'hbf5c61a1;
    ram_cell[     587] = 32'h79f5f7b7;
    ram_cell[     588] = 32'h47991c46;
    ram_cell[     589] = 32'hc973acdb;
    ram_cell[     590] = 32'h9117d70a;
    ram_cell[     591] = 32'hf0b60853;
    ram_cell[     592] = 32'h36a72c4b;
    ram_cell[     593] = 32'h55daae7d;
    ram_cell[     594] = 32'h63dfce8f;
    ram_cell[     595] = 32'hbc256cf6;
    ram_cell[     596] = 32'h1e37362f;
    ram_cell[     597] = 32'h7a37670a;
    ram_cell[     598] = 32'h73cc4f56;
    ram_cell[     599] = 32'h89612337;
    ram_cell[     600] = 32'hf7f0e802;
    ram_cell[     601] = 32'h79856362;
    ram_cell[     602] = 32'ha26a1fa8;
    ram_cell[     603] = 32'h14c25a1c;
    ram_cell[     604] = 32'h2c3ce950;
    ram_cell[     605] = 32'h7c75559f;
    ram_cell[     606] = 32'hbe042099;
    ram_cell[     607] = 32'h88aba1f9;
    ram_cell[     608] = 32'he3a7338b;
    ram_cell[     609] = 32'h28ebce1e;
    ram_cell[     610] = 32'hd97248dd;
    ram_cell[     611] = 32'he32a5a46;
    ram_cell[     612] = 32'hc21c970b;
    ram_cell[     613] = 32'h690bf6e5;
    ram_cell[     614] = 32'h2514ce85;
    ram_cell[     615] = 32'h93dafd16;
    ram_cell[     616] = 32'h19234d23;
    ram_cell[     617] = 32'hb60c3522;
    ram_cell[     618] = 32'hf6ad39fa;
    ram_cell[     619] = 32'h66fc5172;
    ram_cell[     620] = 32'ha9640a3e;
    ram_cell[     621] = 32'hdfade70e;
    ram_cell[     622] = 32'h9600c44f;
    ram_cell[     623] = 32'hf5db2d0d;
    ram_cell[     624] = 32'h8d2e961a;
    ram_cell[     625] = 32'h0782bd76;
    ram_cell[     626] = 32'hc5f6cd23;
    ram_cell[     627] = 32'h4a3a7ea3;
    ram_cell[     628] = 32'hc5d627a7;
    ram_cell[     629] = 32'h0975560e;
    ram_cell[     630] = 32'h6f002ea2;
    ram_cell[     631] = 32'hdf537652;
    ram_cell[     632] = 32'h2e281fdd;
    ram_cell[     633] = 32'h5f27ac6b;
    ram_cell[     634] = 32'h81c05a83;
    ram_cell[     635] = 32'h9c77e605;
    ram_cell[     636] = 32'h33528a14;
    ram_cell[     637] = 32'h9f825720;
    ram_cell[     638] = 32'h19040455;
    ram_cell[     639] = 32'h53cbd3ad;
    ram_cell[     640] = 32'h1d992da5;
    ram_cell[     641] = 32'ha6f8f5cd;
    ram_cell[     642] = 32'h6b18f308;
    ram_cell[     643] = 32'h4304925f;
    ram_cell[     644] = 32'hea60f2e2;
    ram_cell[     645] = 32'h6b82b8aa;
    ram_cell[     646] = 32'ha4095643;
    ram_cell[     647] = 32'h6eadb362;
    ram_cell[     648] = 32'hf6d7b999;
    ram_cell[     649] = 32'h17dcd0b9;
    ram_cell[     650] = 32'h4c833339;
    ram_cell[     651] = 32'h8d89d544;
    ram_cell[     652] = 32'hfb07053d;
    ram_cell[     653] = 32'h35745c46;
    ram_cell[     654] = 32'h392b2164;
    ram_cell[     655] = 32'hd2ff5088;
    ram_cell[     656] = 32'h74760d28;
    ram_cell[     657] = 32'hdc7045e0;
    ram_cell[     658] = 32'h6ac76d25;
    ram_cell[     659] = 32'h078d5d0b;
    ram_cell[     660] = 32'haa4c65c1;
    ram_cell[     661] = 32'h748c3e42;
    ram_cell[     662] = 32'h83bf6d72;
    ram_cell[     663] = 32'hd04c8426;
    ram_cell[     664] = 32'h7f1b6309;
    ram_cell[     665] = 32'h5cc8587f;
    ram_cell[     666] = 32'h2e812ed6;
    ram_cell[     667] = 32'h7457fb19;
    ram_cell[     668] = 32'h0b50dd34;
    ram_cell[     669] = 32'he7fa19a5;
    ram_cell[     670] = 32'hd3867974;
    ram_cell[     671] = 32'he8f4b731;
    ram_cell[     672] = 32'h87733a29;
    ram_cell[     673] = 32'h662fa63e;
    ram_cell[     674] = 32'hecc20aa7;
    ram_cell[     675] = 32'hb3c8d71b;
    ram_cell[     676] = 32'h7ca53bf2;
    ram_cell[     677] = 32'ha3fcb6cf;
    ram_cell[     678] = 32'h8f6f6f2c;
    ram_cell[     679] = 32'h5285f3a1;
    ram_cell[     680] = 32'h765b851d;
    ram_cell[     681] = 32'he443b53e;
    ram_cell[     682] = 32'hc007befd;
    ram_cell[     683] = 32'h9856040e;
    ram_cell[     684] = 32'h52f401f0;
    ram_cell[     685] = 32'hdf0cdf9a;
    ram_cell[     686] = 32'hcf9b15e8;
    ram_cell[     687] = 32'h1c164b9f;
    ram_cell[     688] = 32'hc725eef5;
    ram_cell[     689] = 32'hd34d5884;
    ram_cell[     690] = 32'h85b301d9;
    ram_cell[     691] = 32'h97d1a34a;
    ram_cell[     692] = 32'h70e98bdd;
    ram_cell[     693] = 32'hc1a5c182;
    ram_cell[     694] = 32'ha23ed36d;
    ram_cell[     695] = 32'he4566c2d;
    ram_cell[     696] = 32'hda371f0c;
    ram_cell[     697] = 32'hdbd7968a;
    ram_cell[     698] = 32'he996ccca;
    ram_cell[     699] = 32'hd5429cd6;
    ram_cell[     700] = 32'h30a276c0;
    ram_cell[     701] = 32'hea6782d6;
    ram_cell[     702] = 32'h210c1085;
    ram_cell[     703] = 32'he61e4e2d;
    ram_cell[     704] = 32'h62a62a67;
    ram_cell[     705] = 32'h38f30f29;
    ram_cell[     706] = 32'he49c82bc;
    ram_cell[     707] = 32'h16cec9fc;
    ram_cell[     708] = 32'h00e588e5;
    ram_cell[     709] = 32'h850da34f;
    ram_cell[     710] = 32'h86374365;
    ram_cell[     711] = 32'hd8ba804c;
    ram_cell[     712] = 32'hd5474612;
    ram_cell[     713] = 32'hf08b7a5d;
    ram_cell[     714] = 32'hd1c26bca;
    ram_cell[     715] = 32'h2c32cc70;
    ram_cell[     716] = 32'h619420c3;
    ram_cell[     717] = 32'h45628fbb;
    ram_cell[     718] = 32'hbe60c266;
    ram_cell[     719] = 32'h93f28120;
    ram_cell[     720] = 32'hda3a37d1;
    ram_cell[     721] = 32'hfa8991ec;
    ram_cell[     722] = 32'h7dfe3975;
    ram_cell[     723] = 32'h2524df29;
    ram_cell[     724] = 32'hbb1503ce;
    ram_cell[     725] = 32'hd680ba4f;
    ram_cell[     726] = 32'he7e13d8a;
    ram_cell[     727] = 32'h4782bec9;
    ram_cell[     728] = 32'h326bef46;
    ram_cell[     729] = 32'h3c4adf07;
    ram_cell[     730] = 32'h32dc146d;
    ram_cell[     731] = 32'h051f4695;
    ram_cell[     732] = 32'ha6280b35;
    ram_cell[     733] = 32'h5c2a1150;
    ram_cell[     734] = 32'h0b151596;
    ram_cell[     735] = 32'h3c471cc8;
    ram_cell[     736] = 32'he02badee;
    ram_cell[     737] = 32'h2f985c6d;
    ram_cell[     738] = 32'hec2eedf5;
    ram_cell[     739] = 32'h1a02a2da;
    ram_cell[     740] = 32'h46ca4fb3;
    ram_cell[     741] = 32'hd39e7c12;
    ram_cell[     742] = 32'h8912fbca;
    ram_cell[     743] = 32'he868d823;
    ram_cell[     744] = 32'h72e8a66d;
    ram_cell[     745] = 32'h431f0a94;
    ram_cell[     746] = 32'h7e3225d7;
    ram_cell[     747] = 32'h0b409ae2;
    ram_cell[     748] = 32'h8e976234;
    ram_cell[     749] = 32'h43af991e;
    ram_cell[     750] = 32'h3836dab2;
    ram_cell[     751] = 32'h6c5f3951;
    ram_cell[     752] = 32'h997cd0f6;
    ram_cell[     753] = 32'ha0a75b62;
    ram_cell[     754] = 32'h2b42675d;
    ram_cell[     755] = 32'he0efa570;
    ram_cell[     756] = 32'h8250a04e;
    ram_cell[     757] = 32'h23acff0a;
    ram_cell[     758] = 32'he2df7a9c;
    ram_cell[     759] = 32'h331e6b97;
    ram_cell[     760] = 32'hcb4ff38f;
    ram_cell[     761] = 32'hf2e1134e;
    ram_cell[     762] = 32'ha75b8185;
    ram_cell[     763] = 32'he5e25b42;
    ram_cell[     764] = 32'h8377673c;
    ram_cell[     765] = 32'haea59796;
    ram_cell[     766] = 32'hbeed0ea5;
    ram_cell[     767] = 32'h9139bf3c;
end

endmodule

